library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testcircuit_test is
end testcircuit_test;

architecture test of testcircuit_test is

component TestCircuit
generic (
         Nbit: Integer := 8;
         Mbit: Natural := 16);
port (
      IN1: IN std_logic_vector(Nbit-1 downto 0);
      IN2: IN std_logic_vector(Nbit downto 0);
      IN3: IN std_logic_vector(6 downto 0);
      SEL1: IN std_logic;
      OUT1: OUT std_logic_vector(Mbit-1 downto 0);
      OUT2: OUT std_logic);
end component;

signal IN1_i: std_logic_vector(15 downto 0) := (others => '0');
signal IN2_i: std_logic_vector(16 downto 0) := (others => '0');
signal IN3_i: std_logic_vector(6 downto 0) := (others => '0');
signal SEL1_i: std_logic:= '0';
signal OUT1_i: std_logic_vector(31 downto 0) := (others => '0');
signal OUT2_i: std_logic:= '0';

begin

DUT:TestCircuit
generic map (
             Nbit => 16,
             Mbit => 32)
port map (
          IN1 => IN1_i,
          IN2 => IN2_i,
          IN3 => IN3_i,
          SEL1 => SEL1_i,
          OUT1 => OUT1_i,
          OUT2 => OUT2_i);

TEST: process 

begin 

   IN1_i <= "0110011100010011";
   IN2_i <= "01001111001110010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001110110";
   IN2_i <= "00110000000010110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010011000";
   IN2_i <= "01011001101010101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110101010";
   IN2_i <= "00011011111000111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000001110";
   IN2_i <= "01111100011110110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001111111";
   IN2_i <= "01110110010001111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011101000";
   IN2_i <= "01010100100100000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110101001";
   IN2_i <= "01111111101101010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101000101";
   IN2_i <= "01000010111101100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000111";
   IN2_i <= "01011011101000101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010100100";
   IN2_i <= "01100100010011011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010111001";
   IN2_i <= "00101010100111001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011101001";
   IN2_i <= "00100000100101001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010110010";
   IN2_i <= "00011110011111101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010000001";
   IN2_i <= "01010110001111011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111111000";
   IN2_i <= "00110101101000100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010001101";
   IN2_i <= "01101011010001011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011010110";
   IN2_i <= "01010110010110111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100011011";
   IN2_i <= "00000110100010001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110001110";
   IN2_i <= "00110011111000010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111001000";
   IN2_i <= "00101001100110001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011000100";
   IN2_i <= "00001001011111100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010010110";
   IN2_i <= "01001101001000011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111111";
   IN2_i <= "00001000011110011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100101111";
   IN2_i <= "01000101001100100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110111001";
   IN2_i <= "00010001011010110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010110011";
   IN2_i <= "00101011111000111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000001010";
   IN2_i <= "01000110010110001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101110111";
   IN2_i <= "00100011111011110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000110111";
   IN2_i <= "01011110010011011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010101110";
   IN2_i <= "00111100100000000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001111000";
   IN2_i <= "00000101110111100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110001111";
   IN2_i <= "00011100001101110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100111111";
   IN2_i <= "00110100010011100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111001100";
   IN2_i <= "00100011111001011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101011101";
   IN2_i <= "01000010100001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011111";
   IN2_i <= "01101011010000111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000111011";
   IN2_i <= "01001111001001001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111101011";
   IN2_i <= "00000000010110000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010000110";
   IN2_i <= "01110100111011010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000110000";
   IN2_i <= "00011001010100011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110111110";
   IN2_i <= "01101101010110000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011100010";
   IN2_i <= "00010000001011101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010010001";
   IN2_i <= "00101010001001010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001000111";
   IN2_i <= "01000111010001000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100110101";
   IN2_i <= "00100011011110111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001101100";
   IN2_i <= "01000010111111110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001100010";
   IN2_i <= "01110111001100110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101101101";
   IN2_i <= "01011100011110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110010100";
   IN2_i <= "00010010011010111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010100110";
   IN2_i <= "00001111010010010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101110110";
   IN2_i <= "01010011101101111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111110000";
   IN2_i <= "01010001001000001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001011";
   IN2_i <= "01111011011011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000100";
   IN2_i <= "00010011101110100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100111001";
   IN2_i <= "00011000100100011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011011100";
   IN2_i <= "00010011001110001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011000111";
   IN2_i <= "00010100111000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001011101";
   IN2_i <= "00011000010000010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001010010";
   IN2_i <= "00010001110101001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001101010";
   IN2_i <= "00000110101111011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011101111";
   IN2_i <= "01111100001100011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001010100";
   IN2_i <= "01100111111101101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111000110";
   IN2_i <= "01110001000110011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011011111";
   IN2_i <= "01000001100000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100000010";
   IN2_i <= "01111110010110111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101100010";
   IN2_i <= "00110100001010001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000000101";
   IN2_i <= "00101010110100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111011001";
   IN2_i <= "01011010101001111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011111";
   IN2_i <= "00101111110111010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010010001";
   IN2_i <= "01111011011001111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101101";
   IN2_i <= "01101101100000101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011001110";
   IN2_i <= "01111001111110110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111100011";
   IN2_i <= "00110101001101111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000101010";
   IN2_i <= "01111010100011010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010000100";
   IN2_i <= "01000110000100100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100000";
   IN2_i <= "00011100110010100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100010111";
   IN2_i <= "00111011010010111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011010000";
   IN2_i <= "01000100000110011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100111111";
   IN2_i <= "01100100000101100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011011111";
   IN2_i <= "00000100101101010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010001110";
   IN2_i <= "01000111101000011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101011001";
   IN2_i <= "01010011100000101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100100";
   IN2_i <= "00101101000101010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100101111";
   IN2_i <= "00000010010010100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111100000";
   IN2_i <= "01100000100001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110111001";
   IN2_i <= "00111110101101000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101000011";
   IN2_i <= "00101100111110000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011100001";
   IN2_i <= "01111001010010000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111110001";
   IN2_i <= "01100011001111111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011110011";
   IN2_i <= "00001110110100110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000111111";
   IN2_i <= "00011111101011101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110011011";
   IN2_i <= "01011110110110101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110100101";
   IN2_i <= "00011101001100010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011001001";
   IN2_i <= "01001111111111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110011010";
   IN2_i <= "00101000101101010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101111011";
   IN2_i <= "01001101111011110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110011101";
   IN2_i <= "01000011001111110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101100100";
   IN2_i <= "01111001100011010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100001000";
   IN2_i <= "01011000101010101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101110011";
   IN2_i <= "00110001011111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101111011";
   IN2_i <= "01101100110101111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101100101";
   IN2_i <= "00000000010000000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011110001";
   IN2_i <= "00100100100011000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101001001";
   IN2_i <= "01001111001001100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111110000";
   IN2_i <= "01010110010111101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101111101";
   IN2_i <= "01010010100011001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111100011";
   IN2_i <= "00001001010000100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010010011";
   IN2_i <= "00001010111100000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101011010";
   IN2_i <= "00000010000000110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011111";
   IN2_i <= "00010111101110111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000010001";
   IN2_i <= "00101001001010101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000010";
   IN2_i <= "01010000010101010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011100110";
   IN2_i <= "00100011000101101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010011001";
   IN2_i <= "01001001001010110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000100000";
   IN2_i <= "01011000001010000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101100111";
   IN2_i <= "01011100011010011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010110101";
   IN2_i <= "01111001101000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011100001";
   IN2_i <= "01111001101010011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001001";
   IN2_i <= "00010001000001101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000010011";
   IN2_i <= "00110110011111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011100111";
   IN2_i <= "00001010101111010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000011111";
   IN2_i <= "00110001011010111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101101100";
   IN2_i <= "01000100000010111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101101";
   IN2_i <= "01101110010110011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100110011";
   IN2_i <= "00110010101011100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111110000";
   IN2_i <= "01111101001001001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010010110";
   IN2_i <= "00110100100010000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010010100";
   IN2_i <= "00101110110000100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111000";
   IN2_i <= "01100101010101001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011000100";
   IN2_i <= "00000101000000010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100011000";
   IN2_i <= "01101111000001001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110000111";
   IN2_i <= "00000010101011000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011101110";
   IN2_i <= "00000011001010111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010110";
   IN2_i <= "00001010000110100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001010111";
   IN2_i <= "01101000111011101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000001100";
   IN2_i <= "00011111001111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000101101";
   IN2_i <= "00101101011100001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111111101";
   IN2_i <= "00101100010101010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100100101";
   IN2_i <= "00111011110000101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101111101";
   IN2_i <= "01000010000101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001100111";
   IN2_i <= "01011000100001001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001001111";
   IN2_i <= "00100010011110100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011000011";
   IN2_i <= "01110100111010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001100";
   IN2_i <= "01010001100111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101100010";
   IN2_i <= "00100011010101101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010011";
   IN2_i <= "00110010010111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111110011";
   IN2_i <= "00001011111110111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001111011";
   IN2_i <= "01100111010100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010000101";
   IN2_i <= "00101111000111001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001010001";
   IN2_i <= "01001000111000110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111110110";
   IN2_i <= "01000100001110101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100110001";
   IN2_i <= "00110110010011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100101000";
   IN2_i <= "00100001010001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110011001";
   IN2_i <= "00101111100010011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111001100";
   IN2_i <= "00110101000110101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011001100";
   IN2_i <= "00111010110100001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100011100";
   IN2_i <= "01100011011111100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010101101";
   IN2_i <= "00111010011111011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111111011";
   IN2_i <= "00000010000000110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101001";
   IN2_i <= "00100001101010001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110000011";
   IN2_i <= "01111011001111100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001101001";
   IN2_i <= "00100100111110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011110101";
   IN2_i <= "01111000011100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000101011";
   IN2_i <= "01011111111100000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100000100";
   IN2_i <= "00010010100001001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011011100";
   IN2_i <= "01010000011001100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001110001";
   IN2_i <= "00001110111100011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001110110";
   IN2_i <= "00100011001010110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010100000";
   IN2_i <= "00111100001111101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100111111";
   IN2_i <= "01100110011010011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100011";
   IN2_i <= "01110010111111111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100100100";
   IN2_i <= "00010001100010001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010011111";
   IN2_i <= "00011111111011100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011110";
   IN2_i <= "01010101010101001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110100010";
   IN2_i <= "00000000111000000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000100101";
   IN2_i <= "00101100110101100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101010110";
   IN2_i <= "00001101001101010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111011001";
   IN2_i <= "00001011110001100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001011100";
   IN2_i <= "01011011000100000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011110101";
   IN2_i <= "01100100111100000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111010011";
   IN2_i <= "01001010110000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101101010";
   IN2_i <= "00000110110010000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011000111";
   IN2_i <= "01011111000011101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001100000";
   IN2_i <= "01110100011110101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101000101";
   IN2_i <= "01011110000010100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001101110";
   IN2_i <= "01010010111011010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111001111";
   IN2_i <= "01011010000001001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100001100";
   IN2_i <= "00101111110001101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010111101";
   IN2_i <= "00000100000111001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000011001";
   IN2_i <= "01100111010111001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101110110";
   IN2_i <= "00000111011011100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000100000";
   IN2_i <= "01110110010100100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001000010";
   IN2_i <= "01011100101010010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010101111";
   IN2_i <= "01100101010000000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110011100";
   IN2_i <= "00010000100010001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011010101";
   IN2_i <= "01011111111101101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010101";
   IN2_i <= "01000111110110001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100001111";
   IN2_i <= "00000001100110011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111100000";
   IN2_i <= "01010110111011100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010101101";
   IN2_i <= "00010011010000011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000110101";
   IN2_i <= "00101001000011110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100001011";
   IN2_i <= "01111001010000100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010000101";
   IN2_i <= "01111100000010110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111111110";
   IN2_i <= "01101011011111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000010101";
   IN2_i <= "01101000101001100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101111000";
   IN2_i <= "01101101101110111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100101010";
   IN2_i <= "01001111101100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101101101";
   IN2_i <= "01001000000000111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110011001";
   IN2_i <= "00111101101110001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000000101";
   IN2_i <= "01101010111000000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001001010";
   IN2_i <= "00011100100001000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011000010";
   IN2_i <= "01100101110011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010110010";
   IN2_i <= "00011001011000011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110001111";
   IN2_i <= "00110110011100110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111110";
   IN2_i <= "01110100000001100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000100000";
   IN2_i <= "00010010110000101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111001110";
   IN2_i <= "00001100000101010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000110011";
   IN2_i <= "00111101100000110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010001011";
   IN2_i <= "01101011001111110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011010111";
   IN2_i <= "01101000011100100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011101000";
   IN2_i <= "01010100001101011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100001111";
   IN2_i <= "00001100000010100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101011111";
   IN2_i <= "01110110000001110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001010011";
   IN2_i <= "01100010110101100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100110010";
   IN2_i <= "01111111111001010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110000011";
   IN2_i <= "01001010110111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100100110";
   IN2_i <= "01011100100000101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011011100";
   IN2_i <= "01011101010010111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000111111";
   IN2_i <= "00100011001111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010111001";
   IN2_i <= "00101000111001101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010101011";
   IN2_i <= "01011110101100010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010110000";
   IN2_i <= "01000011010100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110011001";
   IN2_i <= "01011001111100111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100111001";
   IN2_i <= "00100111110111100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000101000";
   IN2_i <= "01010001110111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011011";
   IN2_i <= "01000111000110110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000101011";
   IN2_i <= "00110110100101111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111000011";
   IN2_i <= "00011110011111101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110100111";
   IN2_i <= "00101110111111110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010110011";
   IN2_i <= "00001101001001001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100001100";
   IN2_i <= "01011100111100111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001100000";
   IN2_i <= "01111001111001001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011101101";
   IN2_i <= "01001011110110100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000111001";
   IN2_i <= "00110010010100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111111110";
   IN2_i <= "01100111100000101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000000011";
   IN2_i <= "00001101000010001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100001001";
   IN2_i <= "00010100011111100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100100111";
   IN2_i <= "01001110111101111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100000010";
   IN2_i <= "00101000011101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000001011";
   IN2_i <= "01100100110111010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011010000";
   IN2_i <= "00001011010010110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100000111";
   IN2_i <= "00010011101010001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101110000";
   IN2_i <= "01000111010111110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111001110";
   IN2_i <= "00010110001000000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001001000";
   IN2_i <= "00101000010110000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111111000";
   IN2_i <= "01111111101110100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011010001";
   IN2_i <= "01101110001111010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000000101";
   IN2_i <= "00101101000110000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111000000";
   IN2_i <= "01000010110111000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000010001";
   IN2_i <= "00000111111101001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100101010";
   IN2_i <= "00011001111011100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011111100";
   IN2_i <= "00000110010111100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110100100";
   IN2_i <= "00001001011100100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110111101";
   IN2_i <= "00011111010100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010010";
   IN2_i <= "01110010101101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100001001";
   IN2_i <= "01100011000000101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100101100";
   IN2_i <= "01111001100011000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001110000";
   IN2_i <= "01101100100101001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100101111";
   IN2_i <= "01011111100111111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101110111";
   IN2_i <= "00111101011000000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001110";
   IN2_i <= "00001110111011111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100101011";
   IN2_i <= "01001011000000101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000010100";
   IN2_i <= "00110001001001011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110010111";
   IN2_i <= "01101100011011000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011000";
   IN2_i <= "00011000110011001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111010110";
   IN2_i <= "00111010111110101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010111";
   IN2_i <= "01001010010001111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101100110";
   IN2_i <= "01010010001100010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111010110";
   IN2_i <= "00110011101011100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000011011";
   IN2_i <= "01000010101010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011010101";
   IN2_i <= "01101101111101000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011100101";
   IN2_i <= "00010101001111000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110101100";
   IN2_i <= "00110110111000101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001110000";
   IN2_i <= "00010001001101111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000010111";
   IN2_i <= "01100110011001100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101000011";
   IN2_i <= "00010010100110101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100010010";
   IN2_i <= "01110111100001111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110010010";
   IN2_i <= "01010011100110000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110011010";
   IN2_i <= "00100100010110100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100101010";
   IN2_i <= "01101000111101100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110010001";
   IN2_i <= "00001010000101000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101111001";
   IN2_i <= "01101011010011100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001011000";
   IN2_i <= "00011111100100000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000110100";
   IN2_i <= "01101011101111110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001001001";
   IN2_i <= "00111010111001110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101111100";
   IN2_i <= "00111000010000000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100011011";
   IN2_i <= "00111001101111000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100101";
   IN2_i <= "00111111001101011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000101100";
   IN2_i <= "01110001011110110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110011001";
   IN2_i <= "00110011111101100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111001111";
   IN2_i <= "00101011101011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010000";
   IN2_i <= "00110011001010011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110100010";
   IN2_i <= "00010010110110010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110011";
   IN2_i <= "01011111100010000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111100011";
   IN2_i <= "00100011001000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000001001";
   IN2_i <= "01111101110000110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010010";
   IN2_i <= "00000000110001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010110100";
   IN2_i <= "01110011000000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010111010";
   IN2_i <= "00110100011110100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110110100";
   IN2_i <= "00001010000010011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000010110";
   IN2_i <= "01101010011110011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101111100";
   IN2_i <= "00011000001101101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100011000";
   IN2_i <= "01000111000010010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000101010";
   IN2_i <= "01111011001011100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010100011";
   IN2_i <= "01000111001011001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111000111";
   IN2_i <= "00110111011110001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111110010";
   IN2_i <= "00110100101000101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010101100";
   IN2_i <= "00000111001101011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011110011";
   IN2_i <= "00111001100110111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011011";
   IN2_i <= "00111011110111110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110000";
   IN2_i <= "01101110100110011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101010110";
   IN2_i <= "00101100110111111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110000100";
   IN2_i <= "00000001101001000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000101111";
   IN2_i <= "00111100111100101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110111010";
   IN2_i <= "00001110101000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100110000";
   IN2_i <= "00001110101100010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000010100";
   IN2_i <= "01110111011010110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011110110";
   IN2_i <= "01110000001100010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100001011";
   IN2_i <= "00100011100010101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101000001";
   IN2_i <= "00000111010000011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001001111";
   IN2_i <= "00110010110001000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011110111";
   IN2_i <= "00010100011110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111001010";
   IN2_i <= "00101011001100111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011011110";
   IN2_i <= "00011010010111000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101110111";
   IN2_i <= "01110010010000011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111010100";
   IN2_i <= "00011001111100011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101010000";
   IN2_i <= "01000101110011001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101011011";
   IN2_i <= "01111001010101010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110101000";
   IN2_i <= "00100001011011101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011110";
   IN2_i <= "00010111100001001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100100111";
   IN2_i <= "00111110111011000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000111";
   IN2_i <= "00101011111000010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001000111";
   IN2_i <= "01100010100101100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011110000";
   IN2_i <= "01000011010110111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000110110";
   IN2_i <= "00110111011001000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101010000";
   IN2_i <= "01001000011110111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110000011";
   IN2_i <= "01011010010000111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100011110";
   IN2_i <= "00110010001010111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010001";
   IN2_i <= "01110100101110100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000100011";
   IN2_i <= "00001010010000000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110011101";
   IN2_i <= "01110101111011101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101100010";
   IN2_i <= "01010110010100100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001000";
   IN2_i <= "00101101100101110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111100101";
   IN2_i <= "01000111000001010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111001101";
   IN2_i <= "01010110101101001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011001111";
   IN2_i <= "00110101101010000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100010111";
   IN2_i <= "01110010111100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000100100";
   IN2_i <= "01100100101001101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110111010";
   IN2_i <= "00101101111011000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100111101";
   IN2_i <= "00011001011110101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010001001";
   IN2_i <= "01101001111100111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010100001";
   IN2_i <= "00100010000000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110110111";
   IN2_i <= "00101100111101100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010000000";
   IN2_i <= "01000010010111101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111000110";
   IN2_i <= "00001110110001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011011101";
   IN2_i <= "00101000111110101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001010";
   IN2_i <= "01111011100001111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100110100";
   IN2_i <= "00100000101101010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001101101";
   IN2_i <= "01111010001000110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001011011";
   IN2_i <= "00010010100100101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101000100";
   IN2_i <= "00101111100010001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111011101";
   IN2_i <= "00010010001101100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001111010";
   IN2_i <= "01010101111110110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111101010";
   IN2_i <= "01111111000101001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110101111";
   IN2_i <= "00000010001010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011010000";
   IN2_i <= "01110110110010011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011000110";
   IN2_i <= "00110101111111011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101010001";
   IN2_i <= "00000110001011010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010110";
   IN2_i <= "00110001001011111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100100100";
   IN2_i <= "00000101001011001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101100111";
   IN2_i <= "00000000110110011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110100";
   IN2_i <= "01111101101010110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000101110";
   IN2_i <= "00101100101001001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010010000";
   IN2_i <= "00011101010011010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000010";
   IN2_i <= "01001101110110000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101001010";
   IN2_i <= "00110010111010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011111001";
   IN2_i <= "01111110100111000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101000001";
   IN2_i <= "01111101011110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100101010";
   IN2_i <= "01111010100111010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001010111";
   IN2_i <= "01101110101000011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011011010";
   IN2_i <= "00101110100001000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110000010";
   IN2_i <= "00001001111110101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010111011";
   IN2_i <= "01011001001011011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111011011";
   IN2_i <= "01001110010010101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010011111";
   IN2_i <= "01011101101101001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001101010";
   IN2_i <= "00101110010100000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111100";
   IN2_i <= "00001001001011001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101001111";
   IN2_i <= "01101000001100000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000101110";
   IN2_i <= "01011001110100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011001111";
   IN2_i <= "01110000001000101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110111";
   IN2_i <= "00000000010101011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100100010";
   IN2_i <= "01010000100100000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010111011";
   IN2_i <= "01101001100010001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011110000";
   IN2_i <= "00101011001110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111011000";
   IN2_i <= "01011100001111010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011111100";
   IN2_i <= "01010101011100110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101010011";
   IN2_i <= "01000011001000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000100101";
   IN2_i <= "01010010001101000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010000010";
   IN2_i <= "00011001111110101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110000001";
   IN2_i <= "01010000110000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111010011";
   IN2_i <= "01100101000001110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100101000";
   IN2_i <= "00010001111111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110001001";
   IN2_i <= "00001001011111101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000011000";
   IN2_i <= "01000111100110110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101100000";
   IN2_i <= "00111001110100010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010110000";
   IN2_i <= "01111011110101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001101000";
   IN2_i <= "00110100101101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001100001";
   IN2_i <= "01000001011001111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010110111";
   IN2_i <= "01100100011111010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010011010";
   IN2_i <= "00101001000111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010000";
   IN2_i <= "01110010001110101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011001011";
   IN2_i <= "01100000111101101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101110100";
   IN2_i <= "00110001011000011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010000010";
   IN2_i <= "00000000111100111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001001";
   IN2_i <= "01011101010001111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110000101";
   IN2_i <= "01100101000100000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101010001";
   IN2_i <= "00000011100111101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000100011";
   IN2_i <= "00111100000100110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010001110";
   IN2_i <= "00110001110101100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111111";
   IN2_i <= "00100000111111100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100011011";
   IN2_i <= "01011111000111010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011101011";
   IN2_i <= "01110010000000110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100010";
   IN2_i <= "00100101001101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110010110";
   IN2_i <= "00000110101000100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110101";
   IN2_i <= "00011110110000110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101100111";
   IN2_i <= "00110011111110100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100111000";
   IN2_i <= "01011111001010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100111101";
   IN2_i <= "01011001010110101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000110000";
   IN2_i <= "01001001010111001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011110100";
   IN2_i <= "01000101101001000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010110110";
   IN2_i <= "00110000110110101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000011100";
   IN2_i <= "01110111001100110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100101001";
   IN2_i <= "01000000100001011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110100001";
   IN2_i <= "00001001001100111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011100110";
   IN2_i <= "01110110010001111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000010101";
   IN2_i <= "00000100000000101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001000101";
   IN2_i <= "01111100100011100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010001001";
   IN2_i <= "00100010010010000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001101011";
   IN2_i <= "00001101000001100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101100101";
   IN2_i <= "00001010101100011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011010100";
   IN2_i <= "01010100111110100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101011010";
   IN2_i <= "01110110100000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101010100";
   IN2_i <= "00011110000011001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011011111";
   IN2_i <= "01101111110000011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111110010";
   IN2_i <= "01100000101100101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000111011";
   IN2_i <= "00101010010011100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100000010";
   IN2_i <= "01111100000001100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100000";
   IN2_i <= "01001010000010100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101010011";
   IN2_i <= "01010101110011000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101111001";
   IN2_i <= "00010101001011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101110001";
   IN2_i <= "01101010001010001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011110000";
   IN2_i <= "01010100100110010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011010000";
   IN2_i <= "01000011011001111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001000";
   IN2_i <= "00010111110101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110001110";
   IN2_i <= "00000000010000000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111000010";
   IN2_i <= "01001000011101110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100010011";
   IN2_i <= "01010011110100001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010001100";
   IN2_i <= "00011000000110100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010011011";
   IN2_i <= "01000000011000110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100100110";
   IN2_i <= "01111101101010010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100110000";
   IN2_i <= "01011111111111001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010100110";
   IN2_i <= "00111110000011110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100100001";
   IN2_i <= "00011101010000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100110011";
   IN2_i <= "00011111001000111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011111";
   IN2_i <= "00010100110111111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110011011";
   IN2_i <= "00100010100101101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111101100";
   IN2_i <= "00110010001110010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001100110";
   IN2_i <= "01110111111000001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100010111";
   IN2_i <= "01111000110111010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010000101";
   IN2_i <= "00101111001111011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100001011";
   IN2_i <= "00000111000000000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000010100";
   IN2_i <= "01010000101100001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110100001";
   IN2_i <= "00111010100111001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000011110";
   IN2_i <= "01101110000010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011011001";
   IN2_i <= "00000101000110000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100011101";
   IN2_i <= "00111110111110100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011011000";
   IN2_i <= "00010011101001110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111011111";
   IN2_i <= "00110001110110011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000010111";
   IN2_i <= "01001010011111110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001000001";
   IN2_i <= "01111101011110000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010101";
   IN2_i <= "01101010000011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101001111";
   IN2_i <= "00001101001101010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100010001";
   IN2_i <= "00101110011010100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101101101";
   IN2_i <= "00001101011000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011101111";
   IN2_i <= "00100101010100000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101101101";
   IN2_i <= "00011111001010000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000100111";
   IN2_i <= "01101100101111110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010111010";
   IN2_i <= "00011110010110000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101000000";
   IN2_i <= "00101111101000000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001111110";
   IN2_i <= "00110101111011110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111011011";
   IN2_i <= "01100011111101101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000110000";
   IN2_i <= "01010101101100100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111100110";
   IN2_i <= "00000100000110001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011110101";
   IN2_i <= "01011001010110011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010100001";
   IN2_i <= "01111100111010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100100110";
   IN2_i <= "00011100011110011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101001111";
   IN2_i <= "00100000001110101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111111111";
   IN2_i <= "00011100101111101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101111011";
   IN2_i <= "00110001110110101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010000";
   IN2_i <= "00010011101010101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001101101";
   IN2_i <= "00011001001111111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110111110";
   IN2_i <= "00010111101011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001011100";
   IN2_i <= "01000110111011111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100000011";
   IN2_i <= "01100110101000100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011010110";
   IN2_i <= "00101110100100011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111101100";
   IN2_i <= "01101100101010000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010001110";
   IN2_i <= "00011111000010100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100000001";
   IN2_i <= "00011101111100100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010001000";
   IN2_i <= "00101110011110001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100111000";
   IN2_i <= "01000111000000001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110001010";
   IN2_i <= "01001110100100011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011011000";
   IN2_i <= "00110011010110010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011100111";
   IN2_i <= "00100001111111011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011000111";
   IN2_i <= "00111011010000000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111110110";
   IN2_i <= "00111011001010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000011";
   IN2_i <= "01101101000111101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011011011";
   IN2_i <= "00110001111010001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111010100";
   IN2_i <= "01111100101111110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010111010";
   IN2_i <= "01001111100100011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100100100";
   IN2_i <= "01100110001101010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000100001";
   IN2_i <= "01101100101101100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010110101";
   IN2_i <= "00101111010011000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011011111";
   IN2_i <= "00111001000011001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010110001";
   IN2_i <= "01001100100010011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011100110";
   IN2_i <= "01001000000000011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111001110";
   IN2_i <= "01001111000010100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000001000";
   IN2_i <= "01111110010101001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001101011";
   IN2_i <= "00100110110111011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011110100";
   IN2_i <= "01000000011101111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110001011";
   IN2_i <= "01011100000001110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110001011";
   IN2_i <= "00000111101001101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011110001";
   IN2_i <= "01010001000010011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110101";
   IN2_i <= "01000010011110111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001110010";
   IN2_i <= "01011000011000100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011111110";
   IN2_i <= "01111110010100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001000110";
   IN2_i <= "00110000010010000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010000111";
   IN2_i <= "01110010111111000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101100000";
   IN2_i <= "00000110101000000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101100110";
   IN2_i <= "00011111001110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100011";
   IN2_i <= "01010001011011101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010001010";
   IN2_i <= "01001101010010011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000000";
   IN2_i <= "01001111011101110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010000100";
   IN2_i <= "01011001000110110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111100100";
   IN2_i <= "00111110000110010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110101110";
   IN2_i <= "00001110111001011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100011011";
   IN2_i <= "00000001011001100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101001101";
   IN2_i <= "00110111111110110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011110101";
   IN2_i <= "01100111101110111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010101001";
   IN2_i <= "00101110111001110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001011010";
   IN2_i <= "00111001101100111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001111";
   IN2_i <= "01001000101101010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010001111";
   IN2_i <= "01100001110001011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101000011";
   IN2_i <= "00011011000011101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110011100";
   IN2_i <= "01001001001010100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101111011";
   IN2_i <= "01010100111011010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101001010";
   IN2_i <= "01100100011010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001100001";
   IN2_i <= "00011000111110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000110100";
   IN2_i <= "01110110001001001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010111011";
   IN2_i <= "01000011001111011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010100100";
   IN2_i <= "00010111011110010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011011110";
   IN2_i <= "00110011010110101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101011001";
   IN2_i <= "00100111101111110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011100101";
   IN2_i <= "01000110010100001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001100010";
   IN2_i <= "00111111110011011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001010000";
   IN2_i <= "00111111011110110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000101111";
   IN2_i <= "00111000011010111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111001011";
   IN2_i <= "01110101111001011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100110111";
   IN2_i <= "01011000011001110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010001100";
   IN2_i <= "00111100111110110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110100101";
   IN2_i <= "00100101010010001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101010000";
   IN2_i <= "01001000100110011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100100010";
   IN2_i <= "01010110111110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110111110";
   IN2_i <= "00000100101001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100000100";
   IN2_i <= "00111101100011110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010011110";
   IN2_i <= "01010011010011100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101011";
   IN2_i <= "00110100000110000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011111000";
   IN2_i <= "01001001001010101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011001000";
   IN2_i <= "00011001110110101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110000000";
   IN2_i <= "01011111100110101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001101100";
   IN2_i <= "01001110100011110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111010001";
   IN2_i <= "01110110111011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010110110";
   IN2_i <= "00010101001110101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110111110";
   IN2_i <= "01011111001010110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011111000";
   IN2_i <= "01100000000100011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000011100";
   IN2_i <= "00100011000100011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101111100";
   IN2_i <= "01011110011001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010001110";
   IN2_i <= "00010001100001010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100111101";
   IN2_i <= "01001111111001000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100111111";
   IN2_i <= "00100111101001001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000110010";
   IN2_i <= "01100011110100101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001100000";
   IN2_i <= "01011001010011011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111110001";
   IN2_i <= "01110100100101010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001100001";
   IN2_i <= "00100110000010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100101011";
   IN2_i <= "01000111101000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110001111";
   IN2_i <= "00111111011011010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100010110";
   IN2_i <= "00101000001010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111011001";
   IN2_i <= "01011100111111100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010110111";
   IN2_i <= "01101111000001100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110110";
   IN2_i <= "00001111001001010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110000111";
   IN2_i <= "01011001111110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110101000";
   IN2_i <= "01011101111101000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111111001";
   IN2_i <= "01101111011110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110111001";
   IN2_i <= "00000011011011110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010011";
   IN2_i <= "01000000100101001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110110100";
   IN2_i <= "00010000111110010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110111000";
   IN2_i <= "00011111000110101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111100101";
   IN2_i <= "00010011111000010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110101100";
   IN2_i <= "00000001011110000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011010110";
   IN2_i <= "00100010001001011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100001010";
   IN2_i <= "00100001010011001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111101";
   IN2_i <= "01010101111000010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010110101";
   IN2_i <= "00111110001010110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110010001";
   IN2_i <= "01110111001111000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010100";
   IN2_i <= "01000100001110011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111111000";
   IN2_i <= "01011010101110000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011100000";
   IN2_i <= "00100000000010110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101101001";
   IN2_i <= "00111011001101001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100010000";
   IN2_i <= "00001111100010001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011110011";
   IN2_i <= "01101010010011011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010010101";
   IN2_i <= "01000110110000101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011001010";
   IN2_i <= "01000000000101010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110111000";
   IN2_i <= "00100000010001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010011100";
   IN2_i <= "00000011110101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100111111";
   IN2_i <= "00000111001100111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110110001";
   IN2_i <= "00100001000000110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111001011";
   IN2_i <= "00101010000000000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111101011";
   IN2_i <= "01010000001110100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110001000";
   IN2_i <= "00000010110011010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000010101";
   IN2_i <= "01011101010011010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001001111";
   IN2_i <= "00111000000011101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011000000";
   IN2_i <= "01000000011100111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010101";
   IN2_i <= "00001111101110010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001100111";
   IN2_i <= "01110100101101001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011000000";
   IN2_i <= "00110000000010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011100110";
   IN2_i <= "01111000000111111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000011011";
   IN2_i <= "01111101101000011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000011100";
   IN2_i <= "01000011100111000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111110111";
   IN2_i <= "00011011011101110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000011110";
   IN2_i <= "01110110011111001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110010100";
   IN2_i <= "00001100010100100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101111";
   IN2_i <= "00000010111110000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001001100";
   IN2_i <= "00010100111101110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100101000";
   IN2_i <= "00101000111100010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111010101";
   IN2_i <= "01110001001001110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000010000";
   IN2_i <= "01010100000000001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101001001";
   IN2_i <= "01000001101000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000001010";
   IN2_i <= "01001011011001100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111001";
   IN2_i <= "01100011000110001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100111011";
   IN2_i <= "00010111100000001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000110000";
   IN2_i <= "01110110011100011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000110110";
   IN2_i <= "01010101101100010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110000001";
   IN2_i <= "00011111001000001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011001011";
   IN2_i <= "00011111101011010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101000111";
   IN2_i <= "00111001101011010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100100111";
   IN2_i <= "00001011000110010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000100011";
   IN2_i <= "01110011000011001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100110100";
   IN2_i <= "00111110000011110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000111101";
   IN2_i <= "00010000011001011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110100000";
   IN2_i <= "01100011110011010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010000110";
   IN2_i <= "01000010101110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110001100";
   IN2_i <= "01101101010110110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101001";
   IN2_i <= "00101001011110010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010110001";
   IN2_i <= "01000100000011101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100000011";
   IN2_i <= "01110000110000011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111111110";
   IN2_i <= "01100001111110111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101000110";
   IN2_i <= "01010010111110101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110100110";
   IN2_i <= "01011000100100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010001";
   IN2_i <= "01101101101100000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000111000";
   IN2_i <= "01111111100010011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110001101";
   IN2_i <= "01001000001111010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101110111";
   IN2_i <= "00111100111001110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100001000";
   IN2_i <= "00100100011110011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101011100";
   IN2_i <= "00000101101010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000010001";
   IN2_i <= "00100110100111010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100101";
   IN2_i <= "00000110110000001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110000101";
   IN2_i <= "00111110010100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100111110";
   IN2_i <= "01111010000111101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011110110";
   IN2_i <= "01110110000000011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111001111";
   IN2_i <= "01010001110110100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011010";
   IN2_i <= "00111011011111001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000101";
   IN2_i <= "01100110100011101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101000000";
   IN2_i <= "00000011100100000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100000011";
   IN2_i <= "00011110111001111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010110101";
   IN2_i <= "00110111101011010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100101001";
   IN2_i <= "01100000011111011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011100";
   IN2_i <= "00001100100111110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101011";
   IN2_i <= "00011100110100001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111100011";
   IN2_i <= "00000101000100011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000111100";
   IN2_i <= "00101110111011010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001001110";
   IN2_i <= "00001111111000110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101101001";
   IN2_i <= "00000000100101010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110000110";
   IN2_i <= "00011110010101110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011011101";
   IN2_i <= "01111110100110110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110010011";
   IN2_i <= "00101111010001011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011111000";
   IN2_i <= "01111111101111000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001011101";
   IN2_i <= "01011001011000100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111100001";
   IN2_i <= "00011101000111100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010011000";
   IN2_i <= "01000001100010011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111100011";
   IN2_i <= "01001010001111001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001100010";
   IN2_i <= "01111101001111010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011110001";
   IN2_i <= "00101010011100110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111000000";
   IN2_i <= "00101100110111110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010101011";
   IN2_i <= "01010100100100111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001011000";
   IN2_i <= "00101000111011111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000110001";
   IN2_i <= "00011101000100101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010110010";
   IN2_i <= "00111000101000101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001010111";
   IN2_i <= "00110000011001000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101110001";
   IN2_i <= "01011010011110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110101001";
   IN2_i <= "00110010011011100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111100010";
   IN2_i <= "00101001000110010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001011100";
   IN2_i <= "00101011100011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010100";
   IN2_i <= "00001110100001110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010101101";
   IN2_i <= "01001010101001010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010101001";
   IN2_i <= "00110111100111100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000101011";
   IN2_i <= "00100101010010100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100110101";
   IN2_i <= "01000110110100101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001101111";
   IN2_i <= "00111000010101011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101001101";
   IN2_i <= "00101001100111011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110011";
   IN2_i <= "01111110011000100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001111011";
   IN2_i <= "01101101000100001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101011011";
   IN2_i <= "01011001011111111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100011001";
   IN2_i <= "00111000101001000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000001110";
   IN2_i <= "00010011001011010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100111111";
   IN2_i <= "00010110101000100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011100011";
   IN2_i <= "00001000110010100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111110111";
   IN2_i <= "00001011001100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010101110";
   IN2_i <= "01000010100101110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111001000";
   IN2_i <= "01001111010010000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101100100";
   IN2_i <= "00010111101101011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111101101";
   IN2_i <= "00111110000110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011011110";
   IN2_i <= "00001001100000010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001000100";
   IN2_i <= "00011101100101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000001100";
   IN2_i <= "01101010110100000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101001011";
   IN2_i <= "01010100011000100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001000";
   IN2_i <= "00110011011110110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011010";
   IN2_i <= "00011001011111011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111101011";
   IN2_i <= "01111001010110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100101000";
   IN2_i <= "00100001001001111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101011001";
   IN2_i <= "00101101001000000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111010111";
   IN2_i <= "00010000101110100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011110011";
   IN2_i <= "01010110010101010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010011";
   IN2_i <= "00010111110001010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100011000";
   IN2_i <= "01110001011011000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000010111";
   IN2_i <= "01010010111110100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110110100";
   IN2_i <= "00110010110110100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110011010";
   IN2_i <= "00001101100001010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111111";
   IN2_i <= "01000111101111001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111110100";
   IN2_i <= "00101110011100101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001000010";
   IN2_i <= "00110001101100010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100100001";
   IN2_i <= "00100010110101111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100101000";
   IN2_i <= "01101001000001001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110110000";
   IN2_i <= "00111011000000101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101110100";
   IN2_i <= "01111001000101011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001100101";
   IN2_i <= "01101000100011100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100110011";
   IN2_i <= "00110011101001010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100010000";
   IN2_i <= "01010111101011100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001010000";
   IN2_i <= "01000101110110000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000100011";
   IN2_i <= "00111010000110110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000011101";
   IN2_i <= "01010110010110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010111101";
   IN2_i <= "01110110110111010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010111000";
   IN2_i <= "00111000010100110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000101011";
   IN2_i <= "00000100011100111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101001100";
   IN2_i <= "01000101011110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110100111";
   IN2_i <= "00001100111010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111011011";
   IN2_i <= "00110111000011100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111110";
   IN2_i <= "01010100011010110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000011111";
   IN2_i <= "00000110110101010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000111011";
   IN2_i <= "00110001010110001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000101";
   IN2_i <= "01111001001110111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100000101";
   IN2_i <= "00001111010010100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011001000";
   IN2_i <= "01001010010110001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001011111";
   IN2_i <= "00000001101011011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010000";
   IN2_i <= "00110101010000000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011001100";
   IN2_i <= "01101110000110000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000011101";
   IN2_i <= "01100100100000001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010001010";
   IN2_i <= "01100010011011010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001110";
   IN2_i <= "00000110111101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101101000";
   IN2_i <= "00010111101111111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011001011";
   IN2_i <= "00010111100011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111000100";
   IN2_i <= "01001111010011101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011000101";
   IN2_i <= "01101100100001000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100100011";
   IN2_i <= "00011100101110100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011111011";
   IN2_i <= "01100000111101010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100110111";
   IN2_i <= "00000111000001001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000010001";
   IN2_i <= "01101101110100010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011000100";
   IN2_i <= "00100100111111100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111001111";
   IN2_i <= "00010111000010001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101010101";
   IN2_i <= "01100101010111001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110110000";
   IN2_i <= "00101000001000000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111011001";
   IN2_i <= "00000001111100010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100001";
   IN2_i <= "00010000011110101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111010110";
   IN2_i <= "00110101111110001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111011111";
   IN2_i <= "00011101100111111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101010011";
   IN2_i <= "01000111100010010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010001100";
   IN2_i <= "00100100101101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110100100";
   IN2_i <= "00110000011010111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110111";
   IN2_i <= "01100100100110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111100101";
   IN2_i <= "01111010111010000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010110100";
   IN2_i <= "00000010010111000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010011011";
   IN2_i <= "00110101101110111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101111001";
   IN2_i <= "00001000010110101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000111010";
   IN2_i <= "00110101110011011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001000";
   IN2_i <= "00010000001101011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101100011";
   IN2_i <= "01110100101111000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011111011";
   IN2_i <= "00110000001011011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010111100";
   IN2_i <= "00101100100001011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100111101";
   IN2_i <= "00011101111011000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110010010";
   IN2_i <= "00010111100000010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111000000";
   IN2_i <= "01001100010101111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100101101";
   IN2_i <= "00110011011101101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001010110";
   IN2_i <= "00111001111110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000100011";
   IN2_i <= "01011000000010100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001010";
   IN2_i <= "00100110110001111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110111010";
   IN2_i <= "01100100110001100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101100001";
   IN2_i <= "00100010110111111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110010001";
   IN2_i <= "01100010110000100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010000000";
   IN2_i <= "01011011101101011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110100001";
   IN2_i <= "01000010100010011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111000011";
   IN2_i <= "01010111111011111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111011001";
   IN2_i <= "00101111100010000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001011011";
   IN2_i <= "01001101000101001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111111101";
   IN2_i <= "00101111011010000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100010011";
   IN2_i <= "00101011101000000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011000000";
   IN2_i <= "00000100000111110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110100110";
   IN2_i <= "01101111101111001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111111111";
   IN2_i <= "01110000101001001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101111";
   IN2_i <= "00110111011110001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111100";
   IN2_i <= "01011010100010011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101010110";
   IN2_i <= "01010011001010101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110010011";
   IN2_i <= "01001010110100100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010010111";
   IN2_i <= "01000110100011000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101000100";
   IN2_i <= "01000001100111101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101110111";
   IN2_i <= "01101100100110001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010010101";
   IN2_i <= "00010010101100111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110110";
   IN2_i <= "01101101111111111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011010001";
   IN2_i <= "01001011010000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100110000";
   IN2_i <= "01001000001010100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111001000";
   IN2_i <= "01011011000111101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010011000";
   IN2_i <= "01101001010111010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111010111";
   IN2_i <= "00101110100100100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101110011";
   IN2_i <= "00110011010101101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000001110";
   IN2_i <= "00010011101000010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111011110";
   IN2_i <= "01100100010100110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101110000";
   IN2_i <= "00110000101010000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110101010";
   IN2_i <= "00101111011101101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001111100";
   IN2_i <= "01001100100101110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111001111";
   IN2_i <= "01001011011101110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101100";
   IN2_i <= "00101000111110001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010101110";
   IN2_i <= "00011010001001111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101000000";
   IN2_i <= "01011111110101101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101111101";
   IN2_i <= "00001000001000011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011010100";
   IN2_i <= "01010001110101110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101110010";
   IN2_i <= "00000010111010000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011000001";
   IN2_i <= "00000100100001010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010010010";
   IN2_i <= "01111001010010010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011110100";
   IN2_i <= "01100001011000100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001101110";
   IN2_i <= "01010110011000010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100100001";
   IN2_i <= "00000101111111111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010101000";
   IN2_i <= "01010011110111011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100110101";
   IN2_i <= "01111000010010111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100000";
   IN2_i <= "00101001101100111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101011110";
   IN2_i <= "00000101100111001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100001101";
   IN2_i <= "01110001100111000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111011111";
   IN2_i <= "01010100111111111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110001111";
   IN2_i <= "01111010010111110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001110100";
   IN2_i <= "01001100111101011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010010101";
   IN2_i <= "01000011000001011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011011001";
   IN2_i <= "00010011010100110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010111100";
   IN2_i <= "01110111001111010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000100000";
   IN2_i <= "01101111001100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010010001";
   IN2_i <= "01011001001001110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010111111";
   IN2_i <= "00110011000100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111000110";
   IN2_i <= "00000011110110011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110010001";
   IN2_i <= "01011101111100101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101000000";
   IN2_i <= "01100011001011100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110101111";
   IN2_i <= "01110101011011110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110101010";
   IN2_i <= "01110100010110010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000010000";
   IN2_i <= "01111011000101110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100100011";
   IN2_i <= "01110010010101111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011100";
   IN2_i <= "01000011111101110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001001101";
   IN2_i <= "00110100110001101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000101101";
   IN2_i <= "01100100100011011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011001000";
   IN2_i <= "00110101011011011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011010001";
   IN2_i <= "01011100100001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011100010";
   IN2_i <= "00100100000011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110010001";
   IN2_i <= "01100000001001100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110110111";
   IN2_i <= "01111011010000101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000000110";
   IN2_i <= "00110010001001001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100000010";
   IN2_i <= "00100111011001101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011100111";
   IN2_i <= "00001011010011100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111111001";
   IN2_i <= "01011100111010011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110000000";
   IN2_i <= "00001100101011010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110110000";
   IN2_i <= "01001000111000101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100100110";
   IN2_i <= "00100101110101010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100110000";
   IN2_i <= "00111110111110110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011110110";
   IN2_i <= "01101000000011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110110100";
   IN2_i <= "00000111110100010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100001111";
   IN2_i <= "01101111010010010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111100001";
   IN2_i <= "01010100110001010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100001";
   IN2_i <= "00001011111001010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000111110";
   IN2_i <= "01101001111111111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011011011";
   IN2_i <= "01100111111011010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101011101";
   IN2_i <= "00000011001001000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101010001";
   IN2_i <= "01010011000101101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010101";
   IN2_i <= "01110110101010011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111111111";
   IN2_i <= "01010010010101001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001110011";
   IN2_i <= "00110000000011100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110000100";
   IN2_i <= "00001100001101111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011110011";
   IN2_i <= "01100000100111001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101001101";
   IN2_i <= "01001000011001111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010100110";
   IN2_i <= "01110010011010000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111000010";
   IN2_i <= "00100100111101101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101110010";
   IN2_i <= "00001010000101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100111000";
   IN2_i <= "00011100000000100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010101000";
   IN2_i <= "00101110000111011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101111011";
   IN2_i <= "00001000011011101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001011101";
   IN2_i <= "00100001001110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001000010";
   IN2_i <= "01100111011000111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001001001";
   IN2_i <= "01001011001011000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001111011";
   IN2_i <= "01001000100100010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000100110";
   IN2_i <= "00000111011010001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110110";
   IN2_i <= "00000101101110111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010000101";
   IN2_i <= "00010000110001100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001010";
   IN2_i <= "01000100111001111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001100001";
   IN2_i <= "00101100011110111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110110101";
   IN2_i <= "01100001111000100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010110";
   IN2_i <= "01101011011010111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000001000";
   IN2_i <= "00101110010110000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101100000";
   IN2_i <= "00000111001101000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001001000";
   IN2_i <= "01001010011000101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101010011";
   IN2_i <= "00111101101110111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101110111";
   IN2_i <= "00111100101101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110100001";
   IN2_i <= "01001001101100001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111100110";
   IN2_i <= "01110110100111010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111010011";
   IN2_i <= "00110000011010111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110010100";
   IN2_i <= "01101011010001011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011100100";
   IN2_i <= "00101111001110110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101111001";
   IN2_i <= "00100001001000000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010010011";
   IN2_i <= "00000000111101101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001111010";
   IN2_i <= "00111110000010010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110110101";
   IN2_i <= "01111101111011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011100000";
   IN2_i <= "00110000010100010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001101110";
   IN2_i <= "01101001010000100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010001010";
   IN2_i <= "00100100001111100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100101110";
   IN2_i <= "01011010101100011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001110";
   IN2_i <= "00110100101101101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001110";
   IN2_i <= "00010011001101000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000010011";
   IN2_i <= "00100011100111010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110101100";
   IN2_i <= "00001111000100110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111111100";
   IN2_i <= "01000000011110011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111100010";
   IN2_i <= "00101101110100001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001000110";
   IN2_i <= "00010001110011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001101";
   IN2_i <= "01110101010110001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000000000";
   IN2_i <= "00010101001011110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111001100";
   IN2_i <= "00100110101000010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000100001";
   IN2_i <= "00100110101011110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001111110";
   IN2_i <= "01011101010110111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100101010";
   IN2_i <= "01101010011010010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101100010";
   IN2_i <= "00111000010000010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110011010";
   IN2_i <= "01000001100100111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101001100";
   IN2_i <= "00011011000100110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011110000";
   IN2_i <= "00010000000011000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010001100";
   IN2_i <= "01111000111100110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111001111";
   IN2_i <= "00100001111100101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111110001";
   IN2_i <= "00011110101000000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000000001";
   IN2_i <= "01111101011100011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000011011";
   IN2_i <= "00111101000001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001111000";
   IN2_i <= "01100100001001111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111111110";
   IN2_i <= "00101101000011000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000000100";
   IN2_i <= "00110111111111010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100111";
   IN2_i <= "00001100100000111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100111101";
   IN2_i <= "01101011000000110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001101";
   IN2_i <= "01011001111111000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000001000";
   IN2_i <= "01101001101011101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000000101";
   IN2_i <= "00010111000001001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011111110";
   IN2_i <= "00100101111100011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001001111";
   IN2_i <= "00010000000010111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101101100";
   IN2_i <= "00001010000000100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011001011";
   IN2_i <= "00110110011011011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111010101";
   IN2_i <= "01010111110101010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001011001";
   IN2_i <= "01110000100101110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100010101";
   IN2_i <= "00110111011011010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001100011";
   IN2_i <= "01111100101000100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011100000";
   IN2_i <= "00111110111010001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101011001";
   IN2_i <= "01110111000110100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010000101";
   IN2_i <= "01100010101100001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110011";
   IN2_i <= "00011100111001011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111110110";
   IN2_i <= "01011111010010010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111001100";
   IN2_i <= "01000011100100000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101101010";
   IN2_i <= "01111010100111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110001";
   IN2_i <= "01101010000110110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111001010";
   IN2_i <= "01001000001011101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111000";
   IN2_i <= "01111111001000011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101110011";
   IN2_i <= "01001111001001011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111110000";
   IN2_i <= "01000101010011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110101111";
   IN2_i <= "01100000001011101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010001000";
   IN2_i <= "00000011100111110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010100111";
   IN2_i <= "00000100110110011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101111010";
   IN2_i <= "00011100001111000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011001110";
   IN2_i <= "01111011100110110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001000001";
   IN2_i <= "00000101101101100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111111111";
   IN2_i <= "00011001111001111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010001";
   IN2_i <= "01001000110011110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110010100";
   IN2_i <= "00001111011110001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010000110";
   IN2_i <= "00011011010011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110100011";
   IN2_i <= "01000011110100010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110011111";
   IN2_i <= "00101110011110100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010000100";
   IN2_i <= "01001011001000101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000101111";
   IN2_i <= "00010101010101101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111101101";
   IN2_i <= "00111001010110100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010111011";
   IN2_i <= "00010101011111010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000010110";
   IN2_i <= "01110111010001011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001111011";
   IN2_i <= "01101000011011000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010000010";
   IN2_i <= "00100111101011011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111101011";
   IN2_i <= "00001000101001000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100101011";
   IN2_i <= "00111111110110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010000100";
   IN2_i <= "01011100101010010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101010001";
   IN2_i <= "00101001000011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000100110";
   IN2_i <= "00110111001100001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111111010";
   IN2_i <= "00011100010001011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110011000";
   IN2_i <= "00111001001111010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000010011";
   IN2_i <= "00010011110010000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101101010";
   IN2_i <= "00010001111001000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111000011";
   IN2_i <= "00100011001110001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000110010";
   IN2_i <= "01101111100001101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110010100";
   IN2_i <= "01100101010011110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000101001";
   IN2_i <= "01010111011001101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100011011";
   IN2_i <= "01101100000100011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001010001";
   IN2_i <= "01100000000000101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000011";
   IN2_i <= "01001100011011001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010111011";
   IN2_i <= "00010000010000011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101010100";
   IN2_i <= "00010001111001101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100101110";
   IN2_i <= "01110110001000011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111101";
   IN2_i <= "01011110011110001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110111111";
   IN2_i <= "00000110110100001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011111001";
   IN2_i <= "01110111110110010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101011111";
   IN2_i <= "00110011010011111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101000001";
   IN2_i <= "01111111011101001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010011001";
   IN2_i <= "01111000101010000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100001001";
   IN2_i <= "00111001001111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111110010";
   IN2_i <= "01001010101101010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100011100";
   IN2_i <= "00001010101011010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100010001";
   IN2_i <= "01010100000110010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100101";
   IN2_i <= "00011111111111001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110001100";
   IN2_i <= "01101100100010000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101001011";
   IN2_i <= "01100011011010100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100001110";
   IN2_i <= "00000011000011111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000000";
   IN2_i <= "00001000011111010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000001001";
   IN2_i <= "01111000010111011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010011";
   IN2_i <= "00110110111110100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111001100";
   IN2_i <= "01110011111011010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011000";
   IN2_i <= "00100101101001000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100101001";
   IN2_i <= "01000001010110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011110000";
   IN2_i <= "00011100000110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111110010";
   IN2_i <= "00100100010101110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100011101";
   IN2_i <= "00110100110110001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001000110";
   IN2_i <= "01010111000000101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110101011";
   IN2_i <= "01111101000000001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100100";
   IN2_i <= "00111111011010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111111100";
   IN2_i <= "01001010101100011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100100010";
   IN2_i <= "01101001011101111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111101100";
   IN2_i <= "00110010101111110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100010100";
   IN2_i <= "00111010010100111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000010011";
   IN2_i <= "00101100111000010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001010001";
   IN2_i <= "00010111101011101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101010010";
   IN2_i <= "01101011000100110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111110101";
   IN2_i <= "00101111100100101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010000000";
   IN2_i <= "01100110111000110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100001010";
   IN2_i <= "01001010100000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100001001";
   IN2_i <= "00000010110100000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000000100";
   IN2_i <= "00100110001011101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111010000";
   IN2_i <= "00011100011010000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110011011";
   IN2_i <= "01001110111110110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000100001";
   IN2_i <= "01011001101001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110000111";
   IN2_i <= "01010000001111100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001000001";
   IN2_i <= "01000000001001001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001011001";
   IN2_i <= "01000111001000110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100100011";
   IN2_i <= "01111001010111000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001001101";
   IN2_i <= "00000100001011101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000010";
   IN2_i <= "01101001000101110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001001101";
   IN2_i <= "00111110101001001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011100100";
   IN2_i <= "01001110110111011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101100";
   IN2_i <= "01111111011011100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001101111";
   IN2_i <= "00001010001110101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011101100";
   IN2_i <= "01010000110111010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100110010";
   IN2_i <= "01101101101011101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001100101";
   IN2_i <= "00010101101010010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010010110";
   IN2_i <= "00011111011000001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111011011";
   IN2_i <= "01111101000110101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101110100";
   IN2_i <= "01010000000000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010100010";
   IN2_i <= "00000110101110010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100111";
   IN2_i <= "00101100110100010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110011101";
   IN2_i <= "00110011000101010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100110110";
   IN2_i <= "00110001010100100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111001000";
   IN2_i <= "01101000110001011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011101111";
   IN2_i <= "00101000110101010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010001111";
   IN2_i <= "01100001100011011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110111001";
   IN2_i <= "01111011000001010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000011111";
   IN2_i <= "00000010111100101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111111000";
   IN2_i <= "01110001010001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101011111";
   IN2_i <= "00010000100010110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110010";
   IN2_i <= "00001011110010110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101101100";
   IN2_i <= "00101100000100110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010000";
   IN2_i <= "01010100011111101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001111010";
   IN2_i <= "00110101101010011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011110011";
   IN2_i <= "00011111101111011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101011001";
   IN2_i <= "00001100010111000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101011";
   IN2_i <= "00001011001100101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101000001";
   IN2_i <= "00011110110111110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000010001";
   IN2_i <= "01001011101110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101010100";
   IN2_i <= "01010110000000110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101111001";
   IN2_i <= "01101001100100100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000010101";
   IN2_i <= "01010001010100101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100111101";
   IN2_i <= "01010110111110101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001101100";
   IN2_i <= "00100101110101000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001001101";
   IN2_i <= "00111010001001001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100001101";
   IN2_i <= "01100000100101001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101011100";
   IN2_i <= "00101011110111010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101010100";
   IN2_i <= "01001010001100110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010101101";
   IN2_i <= "01110101010010000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011100000";
   IN2_i <= "01011000010100010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011001101";
   IN2_i <= "01010001001010000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011011110";
   IN2_i <= "00110101100001100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100011000";
   IN2_i <= "01011010001111000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010101010";
   IN2_i <= "01001000101111100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101011111";
   IN2_i <= "01101100000111101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111111011";
   IN2_i <= "01010010000011011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010010";
   IN2_i <= "00111110011011001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100110110";
   IN2_i <= "00001110000110100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110101110";
   IN2_i <= "01000000001010110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100000010";
   IN2_i <= "00011000101101111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011001101";
   IN2_i <= "00111110010101000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011110000";
   IN2_i <= "00111010101110111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111011100";
   IN2_i <= "00010011011110111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111011000";
   IN2_i <= "00000110100110111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101001110";
   IN2_i <= "01110000011101101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001101000";
   IN2_i <= "01000111101110000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100101000";
   IN2_i <= "00100011001100101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011111101";
   IN2_i <= "00011100001110000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011110000";
   IN2_i <= "01001100000000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001110";
   IN2_i <= "00100111100010011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111000111";
   IN2_i <= "00010000000010100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001110100";
   IN2_i <= "01001101011101110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101010";
   IN2_i <= "00000001110110111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111010111";
   IN2_i <= "00000011000110010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101100101";
   IN2_i <= "01000011000000010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001111001";
   IN2_i <= "00000000010010101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100100100";
   IN2_i <= "01111111011111100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001001";
   IN2_i <= "01100000101011100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110001000";
   IN2_i <= "00001111101110110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101101";
   IN2_i <= "01110001001110111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010101";
   IN2_i <= "00110101010010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100111111";
   IN2_i <= "01110000101001110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101001111";
   IN2_i <= "01101010011001000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011000010";
   IN2_i <= "01011111101110100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011010100";
   IN2_i <= "01010000001000001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101111111";
   IN2_i <= "00100100011110010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101101111";
   IN2_i <= "00011111100001000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111110001";
   IN2_i <= "00100001010011000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111010101";
   IN2_i <= "01001000101110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011111011";
   IN2_i <= "00001110010001000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011110001";
   IN2_i <= "00100010111111000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100100101";
   IN2_i <= "00101101111010000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010110010";
   IN2_i <= "01000111010010010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110001101";
   IN2_i <= "01100000010100110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010110010";
   IN2_i <= "00011011100100000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101001011";
   IN2_i <= "00011100010011110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110010101";
   IN2_i <= "00110011011111011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001011100";
   IN2_i <= "01010110110101011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101110011";
   IN2_i <= "00001111010110100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010001101";
   IN2_i <= "01000011111010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101101100";
   IN2_i <= "01101110010010100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011010000";
   IN2_i <= "00001100011111101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011011111";
   IN2_i <= "00011000100111101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101111011";
   IN2_i <= "01011001101101100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101000";
   IN2_i <= "01101100010111111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110101010";
   IN2_i <= "01000010111100010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001111010";
   IN2_i <= "00000111111011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010001010";
   IN2_i <= "00001001101001011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101100101";
   IN2_i <= "00110000100011010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110111101";
   IN2_i <= "01000011110010000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011100001";
   IN2_i <= "01101100011101000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111000110";
   IN2_i <= "00100001111110101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111100101";
   IN2_i <= "00100000111011101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010011010";
   IN2_i <= "01011111001100001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000011100";
   IN2_i <= "01101101010010000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001111010";
   IN2_i <= "00111010101111101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010101000";
   IN2_i <= "00000000010100000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011101111";
   IN2_i <= "01011011000010100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010100";
   IN2_i <= "01111110110101001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100101100";
   IN2_i <= "01001001001100101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101001010";
   IN2_i <= "00010100011111100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100010101";
   IN2_i <= "01001010000101010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110110010";
   IN2_i <= "00000100000010001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011100001";
   IN2_i <= "00011101111111000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000110111";
   IN2_i <= "01001101000101011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101010111";
   IN2_i <= "01100110011110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110111011";
   IN2_i <= "00000110000101101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110010111";
   IN2_i <= "01010001100101001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000011000";
   IN2_i <= "01001001111001001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100011001";
   IN2_i <= "00001010000000110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001000111";
   IN2_i <= "01000001000010111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010011100";
   IN2_i <= "01001000010101001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111000110";
   IN2_i <= "00010111100110000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101010010";
   IN2_i <= "00001111001001110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010110111";
   IN2_i <= "01111011011011100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111110101";
   IN2_i <= "01011001110100110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111110000";
   IN2_i <= "01001101011000101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101001001";
   IN2_i <= "01000011010110100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000000110";
   IN2_i <= "01111011011010011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111101000";
   IN2_i <= "00000111111001100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001011011";
   IN2_i <= "00000000011010111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011101101";
   IN2_i <= "01000110110101111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101101010";
   IN2_i <= "01000110011111100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100001000";
   IN2_i <= "00110100100110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001110011";
   IN2_i <= "00001110010101110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110111010";
   IN2_i <= "00100001010110011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100010110";
   IN2_i <= "00101001001100111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111101111";
   IN2_i <= "01001101010000000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110011111";
   IN2_i <= "00000000100100001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011010111";
   IN2_i <= "01111011100110011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000011010";
   IN2_i <= "01001111010011101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001001010";
   IN2_i <= "00000001100110110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011010001";
   IN2_i <= "00100011111000110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001001110";
   IN2_i <= "01000001001111101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011101101";
   IN2_i <= "01111010111111100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110101101";
   IN2_i <= "01100100101000100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000100";
   IN2_i <= "01001101001010100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011010000";
   IN2_i <= "01000101011001000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100000010";
   IN2_i <= "01001000111000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101000";
   IN2_i <= "00011011100001000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110101010";
   IN2_i <= "01101001110111000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010111100";
   IN2_i <= "01010101000000010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100000100";
   IN2_i <= "01111010110001100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000010111";
   IN2_i <= "00010111001111100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110011";
   IN2_i <= "01101000101111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100110101";
   IN2_i <= "01011001111010101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100000000";
   IN2_i <= "00100010110100010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010001100";
   IN2_i <= "00011010110110010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000000100";
   IN2_i <= "01110001001000110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010111110";
   IN2_i <= "01001001100100111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110001101";
   IN2_i <= "00111111010100100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011101111";
   IN2_i <= "00101001001010010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000100110";
   IN2_i <= "00110100010000000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010110010";
   IN2_i <= "01101111011101011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100010110";
   IN2_i <= "00101110000001010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011111100";
   IN2_i <= "00110010011000101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110111010";
   IN2_i <= "01110101000001100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100111111";
   IN2_i <= "00001111101110010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101111010";
   IN2_i <= "01001111001110001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110111";
   IN2_i <= "00000010011111110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111100100";
   IN2_i <= "00111010000111100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001100001";
   IN2_i <= "00001001100001110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000001101";
   IN2_i <= "00111010010010111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010001111";
   IN2_i <= "01001110000000000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010010111";
   IN2_i <= "01110010001110001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100110";
   IN2_i <= "00100110110101000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011110000";
   IN2_i <= "00001000010100010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110110010";
   IN2_i <= "01101111001010111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111001110";
   IN2_i <= "00100111101011001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001110100";
   IN2_i <= "00010001110011110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000111001";
   IN2_i <= "01110011110111000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010000000";
   IN2_i <= "00011111011001010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000100001";
   IN2_i <= "00011110000001111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000111010";
   IN2_i <= "00111100010100111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011101110";
   IN2_i <= "00000010010100001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010111110";
   IN2_i <= "00011011110110001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011110100";
   IN2_i <= "01000110010010111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000011001";
   IN2_i <= "01100011100010011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011010000";
   IN2_i <= "00000101000010000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011011010";
   IN2_i <= "01101110100111111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001110001";
   IN2_i <= "00011011101001010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001100100";
   IN2_i <= "01010110111010000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010101111";
   IN2_i <= "01100010010001010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000001110";
   IN2_i <= "01001001100000111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000001000";
   IN2_i <= "01111100101001101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100111101";
   IN2_i <= "01010011010101000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000110011";
   IN2_i <= "01001011010111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100111001";
   IN2_i <= "00111011101100100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000011000";
   IN2_i <= "01110001000010111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111011000";
   IN2_i <= "01111100011100011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110101000";
   IN2_i <= "01110001101110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111000100";
   IN2_i <= "01110110101110010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001011001";
   IN2_i <= "01101011111110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100101";
   IN2_i <= "01000001011100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100111011";
   IN2_i <= "01110011010010100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011010111";
   IN2_i <= "00100010010011011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011101000";
   IN2_i <= "01101010100101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111101101";
   IN2_i <= "01000000111100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100010111";
   IN2_i <= "01010100000010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111001010";
   IN2_i <= "00111001010011010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000100000";
   IN2_i <= "01010001011101100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011110000";
   IN2_i <= "00100010110010010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000001111";
   IN2_i <= "01010011000011111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001100001";
   IN2_i <= "01011110101101011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100111000";
   IN2_i <= "01001010111111011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010111101";
   IN2_i <= "00101001011011010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011001100";
   IN2_i <= "00001010010100011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111111011";
   IN2_i <= "01010100000001001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010110110";
   IN2_i <= "01110000010011001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101101000";
   IN2_i <= "01110110111101000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011011010";
   IN2_i <= "00110100100011111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100000101";
   IN2_i <= "00100010010001001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100000001";
   IN2_i <= "00100000011100101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111111110";
   IN2_i <= "00101110100111111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010010101";
   IN2_i <= "01011100111101101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010111010";
   IN2_i <= "01010000001111001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110100110";
   IN2_i <= "00011010010011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110110111";
   IN2_i <= "01010100010100111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101001101";
   IN2_i <= "01000010010101010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100100100";
   IN2_i <= "00101001010010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110111";
   IN2_i <= "01110100001010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101011111";
   IN2_i <= "00100011100100101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001110010";
   IN2_i <= "01001011111000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110011001";
   IN2_i <= "01010010010111010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011010010";
   IN2_i <= "01000000010111001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111101100";
   IN2_i <= "00110011001110100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000010111";
   IN2_i <= "00001111111000110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010110001";
   IN2_i <= "01011110111011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011001111";
   IN2_i <= "00101111001010110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110100001";
   IN2_i <= "01010100110100001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101111001";
   IN2_i <= "00111010011010011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101010110";
   IN2_i <= "01011110010001011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111010011";
   IN2_i <= "01011010011111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000001011";
   IN2_i <= "01001011101101001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011110111";
   IN2_i <= "01010111001111000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111101011";
   IN2_i <= "00001010100000001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010010100";
   IN2_i <= "01010111110011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011001011";
   IN2_i <= "00111110010111110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100010011";
   IN2_i <= "01001001100111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011111";
   IN2_i <= "00111111010101110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110011";
   IN2_i <= "00010001010001110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101100011";
   IN2_i <= "00111100011011010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011001100";
   IN2_i <= "00111100101111110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111101010";
   IN2_i <= "00100000000011011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010010101";
   IN2_i <= "01001111010011110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011010110";
   IN2_i <= "01111110111111100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000010010";
   IN2_i <= "00001010011010101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110001110";
   IN2_i <= "01101100011011100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010101111";
   IN2_i <= "01001011101110110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001011010";
   IN2_i <= "01000111010010101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101010010";
   IN2_i <= "00101000000001001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100111";
   IN2_i <= "00000111100110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110100011";
   IN2_i <= "01011001001000001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011000000";
   IN2_i <= "01110011011110100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101101011";
   IN2_i <= "01110001100011111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001000101";
   IN2_i <= "01011001101010001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010001000";
   IN2_i <= "01001000101110100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001000";
   IN2_i <= "01110100101010001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101011001";
   IN2_i <= "00110101011101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101000110";
   IN2_i <= "00111101110111000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000100010";
   IN2_i <= "01010000010011001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111010010";
   IN2_i <= "00100001001110001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110100111";
   IN2_i <= "00100000011111111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000000101";
   IN2_i <= "00011001011010101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110000101";
   IN2_i <= "00100011000010001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010010001";
   IN2_i <= "01100110000110010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000101001";
   IN2_i <= "01001010010010101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111010011";
   IN2_i <= "00001111101000011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100001111";
   IN2_i <= "00110100011101110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100101010";
   IN2_i <= "00001001001100001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010001111";
   IN2_i <= "01100010010100011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101101100";
   IN2_i <= "01001011011111011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110011100";
   IN2_i <= "01001001011000000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011110100";
   IN2_i <= "01100011101101111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011100000";
   IN2_i <= "00011001101011110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000000010";
   IN2_i <= "01001011101111011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110111001";
   IN2_i <= "01001110010010011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000101000";
   IN2_i <= "00000100100101000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110010001";
   IN2_i <= "01100011110011010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111000101";
   IN2_i <= "00110011010010011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010010110";
   IN2_i <= "00101011000010100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111111010";
   IN2_i <= "01010011001101000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000000101";
   IN2_i <= "00110111101100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110101101";
   IN2_i <= "00010010001001100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101111001";
   IN2_i <= "00000010101011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010100111";
   IN2_i <= "00111001110001010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000011001";
   IN2_i <= "01101001101001001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101000000";
   IN2_i <= "01001011111101110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011010110";
   IN2_i <= "00001001111111011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110010101";
   IN2_i <= "01111111001010101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000010001";
   IN2_i <= "01000010100101100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000110101";
   IN2_i <= "00111101000100111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010111101";
   IN2_i <= "00000001100010110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000110100";
   IN2_i <= "01010100010111100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010000000";
   IN2_i <= "01100001100111101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000100010";
   IN2_i <= "01101011111100011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100010011";
   IN2_i <= "00010011110010100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001111011";
   IN2_i <= "00001110111001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001010000";
   IN2_i <= "01100010101110000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010010110";
   IN2_i <= "00000011100000111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100100110";
   IN2_i <= "00100010001111101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101111010";
   IN2_i <= "01100010111101100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110000110";
   IN2_i <= "01011110101110001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110111101";
   IN2_i <= "00100010000011001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001011101";
   IN2_i <= "00101001000100110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011000101";
   IN2_i <= "00101011110010111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010001100";
   IN2_i <= "00110010110110101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000010101";
   IN2_i <= "01001100010000100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111000000";
   IN2_i <= "01010110011000001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111110100";
   IN2_i <= "01100010000011101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111110111";
   IN2_i <= "01000011011001101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111110101";
   IN2_i <= "01011000100111111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111110";
   IN2_i <= "01100101111111101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011101101";
   IN2_i <= "01101110000011100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001011010";
   IN2_i <= "00111001001001100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100100110";
   IN2_i <= "01111001111111010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100101000";
   IN2_i <= "01100011011001000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111001100";
   IN2_i <= "01011011001110011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000010100";
   IN2_i <= "01111111101000011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110111001";
   IN2_i <= "00100111100010010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011101010";
   IN2_i <= "01010101111110000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101011010";
   IN2_i <= "00110000101101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001101000";
   IN2_i <= "00000101010000001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010111111";
   IN2_i <= "00111011000101001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001010";
   IN2_i <= "01101101000010101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010110001";
   IN2_i <= "00000000111101001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001101100";
   IN2_i <= "01011110010000111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000000100";
   IN2_i <= "00000011111101011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100001110";
   IN2_i <= "00110100000000011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111000000";
   IN2_i <= "00010100100100010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101011111";
   IN2_i <= "01011000010011010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101001111";
   IN2_i <= "00001110101110000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100101110";
   IN2_i <= "01000101011000001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110010100";
   IN2_i <= "01011010010010101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000100111";
   IN2_i <= "01001011000101000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100111110";
   IN2_i <= "00011011001010011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100101011";
   IN2_i <= "00001000001111010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000101111";
   IN2_i <= "00001001101110110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000111111";
   IN2_i <= "01100000001000100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001010001";
   IN2_i <= "00110100000110101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010101111";
   IN2_i <= "00111010110001100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101011100";
   IN2_i <= "01000000011000100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001001";
   IN2_i <= "01001000010110100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110011011";
   IN2_i <= "01011000110101010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110010010";
   IN2_i <= "01100110000000001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011001111";
   IN2_i <= "01001111111010010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000100000";
   IN2_i <= "01001111010111110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110110111";
   IN2_i <= "00111100011100011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111011000";
   IN2_i <= "01001111010111000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111110111";
   IN2_i <= "00011101000100000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010101001";
   IN2_i <= "00111010101111101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011010100";
   IN2_i <= "00000011001101110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000110001";
   IN2_i <= "00000110111011010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010011010";
   IN2_i <= "00000000101010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010000011";
   IN2_i <= "01111110010001001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000000101";
   IN2_i <= "01110110000111001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111001101";
   IN2_i <= "01110011110001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110000000";
   IN2_i <= "01010100100001010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101101100";
   IN2_i <= "01111000100010101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010001";
   IN2_i <= "00000011000100111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000110010";
   IN2_i <= "01100000001011101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101001101";
   IN2_i <= "01100001111100111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110011";
   IN2_i <= "01110110001100001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010100011";
   IN2_i <= "00010010001101101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110110011";
   IN2_i <= "01001010100100110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110111110";
   IN2_i <= "01101011001010010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000101101";
   IN2_i <= "00110001100001110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101001100";
   IN2_i <= "01001011011111110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001000000";
   IN2_i <= "01111000101001000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101110010";
   IN2_i <= "00001111000010101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010100000";
   IN2_i <= "00100100011010011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100011";
   IN2_i <= "00110000010001001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000100010";
   IN2_i <= "00010001110111100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111000011";
   IN2_i <= "00011100011110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100101";
   IN2_i <= "01000110100110100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110100100";
   IN2_i <= "00010101110110100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101111001";
   IN2_i <= "01010010111000100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011010001";
   IN2_i <= "00000000101010100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111000110";
   IN2_i <= "00110110001001000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101101110";
   IN2_i <= "00101010011101111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010011110";
   IN2_i <= "01011011111011010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000111000";
   IN2_i <= "01010001111100111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110110100";
   IN2_i <= "00100000010101101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000111100";
   IN2_i <= "01101001111010011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100011011";
   IN2_i <= "01101011101100111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010011110";
   IN2_i <= "01001011111101000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000100001";
   IN2_i <= "00101110000010110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010111110";
   IN2_i <= "00100101101001001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111100001";
   IN2_i <= "01010001100000100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010110000";
   IN2_i <= "00100011101100010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010001000";
   IN2_i <= "00101010000110110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111010010";
   IN2_i <= "01101100111110011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111110010";
   IN2_i <= "01111011000111000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110001111";
   IN2_i <= "00111111110000011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100101110";
   IN2_i <= "00111110010110011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101010111";
   IN2_i <= "00011111101000101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111000";
   IN2_i <= "00111000001010001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011010111";
   IN2_i <= "00001110101000001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011001001";
   IN2_i <= "00011011111100100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101010110";
   IN2_i <= "00010100001111110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111100";
   IN2_i <= "00011010010010111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101111110";
   IN2_i <= "00001101010000110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110011110";
   IN2_i <= "01110000101110001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001000010";
   IN2_i <= "00101010100100001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001100111";
   IN2_i <= "01011110010100011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011011110";
   IN2_i <= "01001010110110100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101000010";
   IN2_i <= "00110011110101110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100100000";
   IN2_i <= "00010100100010010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100101010";
   IN2_i <= "00011000100011010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010001000";
   IN2_i <= "00010110010011110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010000";
   IN2_i <= "01100001010111010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101010111";
   IN2_i <= "01001010111001111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111100011";
   IN2_i <= "00110101110100110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110110010";
   IN2_i <= "01000000100001001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111011000";
   IN2_i <= "00001010101000111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110010011";
   IN2_i <= "00111001101100111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000111010";
   IN2_i <= "01100100001001010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011111010";
   IN2_i <= "01011101000010000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010101";
   IN2_i <= "01010111000101101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110100111";
   IN2_i <= "01100011111110001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111111001";
   IN2_i <= "00110100101100010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101110011";
   IN2_i <= "00010000100011010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101101111";
   IN2_i <= "00100111111100110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010011";
   IN2_i <= "01010010011000000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100111101";
   IN2_i <= "00110010111110111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110100110";
   IN2_i <= "00110000110011111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000000110";
   IN2_i <= "00001110000000111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010001000";
   IN2_i <= "00111110000000000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100101";
   IN2_i <= "01000111101110111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111101110";
   IN2_i <= "01001110010110001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010010101";
   IN2_i <= "00101011101011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011000000";
   IN2_i <= "01010101001000011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010000010";
   IN2_i <= "01110100011001010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100101";
   IN2_i <= "01000011111011110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110110001";
   IN2_i <= "01011100010000001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101110010";
   IN2_i <= "01101100011110100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111110110";
   IN2_i <= "00100111010101010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001110000";
   IN2_i <= "01101011011001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011010110";
   IN2_i <= "01100000000101001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100000101";
   IN2_i <= "00101110101001111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010100101";
   IN2_i <= "01111010011100110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110011010";
   IN2_i <= "01110000100001110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111110110";
   IN2_i <= "01110010100111000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001001001";
   IN2_i <= "01000101110101001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101100100";
   IN2_i <= "01001001001010100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101001";
   IN2_i <= "00101101000011100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001010000";
   IN2_i <= "00010100111110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100010111";
   IN2_i <= "01001000110111110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010010101";
   IN2_i <= "00100111000011111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101110111";
   IN2_i <= "01110001001111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011011101";
   IN2_i <= "00100001111101010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011001100";
   IN2_i <= "01000101100100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101000001";
   IN2_i <= "00101011011111111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010011001";
   IN2_i <= "01010010110001011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001001110";
   IN2_i <= "00110110111101111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111110011";
   IN2_i <= "01101111000011010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111101111";
   IN2_i <= "00111110100011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100001100";
   IN2_i <= "01101000001110000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001110001";
   IN2_i <= "01101100110011010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010011";
   IN2_i <= "01100010101111001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000001110";
   IN2_i <= "00000011010110001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100100001";
   IN2_i <= "01101001101011000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111101";
   IN2_i <= "01001101000101110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001011111";
   IN2_i <= "01100011110111010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011101011";
   IN2_i <= "00010001010101110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011110110";
   IN2_i <= "01010111100011101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110100001";
   IN2_i <= "01101001000110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011111111";
   IN2_i <= "01001101001010101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001000010";
   IN2_i <= "01010111111011010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101101000";
   IN2_i <= "00100010100011100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100111001";
   IN2_i <= "00110110001100110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010011000";
   IN2_i <= "01001111110001101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010000111";
   IN2_i <= "00000001101001100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010010100";
   IN2_i <= "00100101110110000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110011001";
   IN2_i <= "00000001100010101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000111100";
   IN2_i <= "01110110010010000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100011111";
   IN2_i <= "00110001100010100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111100110";
   IN2_i <= "01001110011111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101000010";
   IN2_i <= "00001000011110001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011100000";
   IN2_i <= "00001001101110101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001100001";
   IN2_i <= "01001100011100001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101000001";
   IN2_i <= "01101010010010100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101000011";
   IN2_i <= "00100011010110101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000010000";
   IN2_i <= "01101010111000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011010";
   IN2_i <= "00111011001000110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110110000";
   IN2_i <= "01110101111000010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011111110";
   IN2_i <= "01011101010110001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111111";
   IN2_i <= "01001101001010011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011100100";
   IN2_i <= "01101111001111000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100010111";
   IN2_i <= "00000011000111000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011000010";
   IN2_i <= "00111001100011010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100100";
   IN2_i <= "00100111001100101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001110010";
   IN2_i <= "00100011010100001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101001011";
   IN2_i <= "00110110111100001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010010000";
   IN2_i <= "00111011110110100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101010";
   IN2_i <= "00111110111101101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000100010";
   IN2_i <= "01010100100010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010000";
   IN2_i <= "01001001110000001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110100000";
   IN2_i <= "00000110001000000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000011100";
   IN2_i <= "01110011010110010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011111011";
   IN2_i <= "01111101110110011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111110101";
   IN2_i <= "01010001000000110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000100000";
   IN2_i <= "01100010000011011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111001101";
   IN2_i <= "00111111001101010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110101110";
   IN2_i <= "00001011110010111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101100";
   IN2_i <= "01100000010011001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100001011";
   IN2_i <= "00010011111000110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000101100";
   IN2_i <= "01101010100010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100001111";
   IN2_i <= "00001100111001100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010100101";
   IN2_i <= "00000111100101011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010001111";
   IN2_i <= "01011100010000111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010010101";
   IN2_i <= "01110000010111011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110101000";
   IN2_i <= "00100110101101100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101110111";
   IN2_i <= "01111101100111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111000001";
   IN2_i <= "00101110000111000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110111110";
   IN2_i <= "01000000101101001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000101111";
   IN2_i <= "00001100000011101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110110010";
   IN2_i <= "01101111011100001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010000001";
   IN2_i <= "01001000011101110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110010010";
   IN2_i <= "01101011100100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000010101";
   IN2_i <= "00011110011110010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110011011";
   IN2_i <= "00010111110010001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011110";
   IN2_i <= "01010100000000111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100011011";
   IN2_i <= "01011011000000000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100100010";
   IN2_i <= "00100001011001011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111010000";
   IN2_i <= "01011000000000101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110011001";
   IN2_i <= "00000100101001011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101010000";
   IN2_i <= "00111111110010010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110110010";
   IN2_i <= "01011011100001111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010000101";
   IN2_i <= "01110011100101100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110110001";
   IN2_i <= "00100000010001101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001000101";
   IN2_i <= "00100010001011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010000000";
   IN2_i <= "01100001000101100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001101111";
   IN2_i <= "01011011110101101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011100011";
   IN2_i <= "01100011101000000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011010001";
   IN2_i <= "00111111001100110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111001010";
   IN2_i <= "01001000001111101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011111010";
   IN2_i <= "01100101000110011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111001100";
   IN2_i <= "01010011111110110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011011000";
   IN2_i <= "00011111111111101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100010";
   IN2_i <= "01110011110110000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000010111";
   IN2_i <= "00101101111011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100011";
   IN2_i <= "01101011000101011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110001100";
   IN2_i <= "00001000111000011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011101101";
   IN2_i <= "01010001011101000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100100";
   IN2_i <= "00000111101011101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100111011";
   IN2_i <= "01001010110010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001010000";
   IN2_i <= "00000100001000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001111011";
   IN2_i <= "00000011010111111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100101100";
   IN2_i <= "00100101100000111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010010100";
   IN2_i <= "00101110100101101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010001000";
   IN2_i <= "01010100111000011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111110101";
   IN2_i <= "00010010010110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011010110";
   IN2_i <= "01000100001111010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111111";
   IN2_i <= "01100101010111010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100000111";
   IN2_i <= "01111011001000000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111111100";
   IN2_i <= "01101110110101010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110110101";
   IN2_i <= "01100001000100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110011110";
   IN2_i <= "01100111000110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111100110";
   IN2_i <= "01110000101010010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011000001";
   IN2_i <= "00100001000101100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001100";
   IN2_i <= "01001111001010100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100011";
   IN2_i <= "00101001001001011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100101011";
   IN2_i <= "00101011001010001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110111111";
   IN2_i <= "01100101111111111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011000011";
   IN2_i <= "01100010011100011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010011011";
   IN2_i <= "01000100111010010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001111100";
   IN2_i <= "00111000011011101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110010110";
   IN2_i <= "00010111011110100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111010110";
   IN2_i <= "00000010111111000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111100";
   IN2_i <= "00011011010101011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111000100";
   IN2_i <= "01111110110000010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011001000";
   IN2_i <= "01101000011101110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101110010";
   IN2_i <= "00000110011110011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111000100";
   IN2_i <= "00011001011111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110011011";
   IN2_i <= "00110000101100001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001000001";
   IN2_i <= "00110100001110010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110110001";
   IN2_i <= "01100000111000010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100010001";
   IN2_i <= "01001001001111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001011010";
   IN2_i <= "01101100001010011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011101111";
   IN2_i <= "00110000100100010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000010010";
   IN2_i <= "01100110010000101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110100010";
   IN2_i <= "01001101011000110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110111111";
   IN2_i <= "00111001110100101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010101";
   IN2_i <= "00101101110101101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001010110";
   IN2_i <= "00010011010000000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011110011";
   IN2_i <= "00110011011010000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110011010";
   IN2_i <= "01100011110111011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111000011";
   IN2_i <= "00111101110101101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110010011";
   IN2_i <= "00010011010100110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101100010";
   IN2_i <= "01111101100011101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110101111";
   IN2_i <= "00101111110110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111010010";
   IN2_i <= "01101010011111011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011011000";
   IN2_i <= "01010011100100101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111111011";
   IN2_i <= "01110000110010001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001110001";
   IN2_i <= "00111001010011100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001110110";
   IN2_i <= "01011101000101101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111111000";
   IN2_i <= "01001011001001110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000100";
   IN2_i <= "00100100101101110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101110110";
   IN2_i <= "00110010010010001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111111110";
   IN2_i <= "00101010100000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001010110";
   IN2_i <= "00100011000001011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101001001";
   IN2_i <= "00111100100011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011011011";
   IN2_i <= "00011111101011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101111111";
   IN2_i <= "01100100001111100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010100011";
   IN2_i <= "00000101010010001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101111111";
   IN2_i <= "00011100011011010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110010000";
   IN2_i <= "00111110101100110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101000110";
   IN2_i <= "00011000010011000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000010";
   IN2_i <= "00111011100011001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000100011";
   IN2_i <= "00010111010101001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010010111";
   IN2_i <= "00001011100101001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001100";
   IN2_i <= "01000001011100110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111111000";
   IN2_i <= "00010111000010111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001001100";
   IN2_i <= "00101000011010011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011110100";
   IN2_i <= "00111111100110100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110010110";
   IN2_i <= "01100100001011100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001110";
   IN2_i <= "00001000001000011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010100011";
   IN2_i <= "00111010000011100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010000010";
   IN2_i <= "00001111000000111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111101010";
   IN2_i <= "00001011100000011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100111111";
   IN2_i <= "00101110111011000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010010";
   IN2_i <= "01110000101101111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001110101";
   IN2_i <= "00110011111101010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110001011";
   IN2_i <= "01100000111010011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010110";
   IN2_i <= "01101101011101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100001";
   IN2_i <= "01110011010000000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101111001";
   IN2_i <= "01101011001001110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110101100";
   IN2_i <= "01011101001100010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110100101";
   IN2_i <= "00000110011110000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101101110";
   IN2_i <= "00000001010011110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010011010";
   IN2_i <= "00011101000100100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000100100";
   IN2_i <= "01001011010101111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001100011";
   IN2_i <= "00100001000101110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010001000";
   IN2_i <= "00011100101100111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000010000";
   IN2_i <= "00111001011001000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000101110";
   IN2_i <= "01010101011000111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111111";
   IN2_i <= "00110000001100100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000000010";
   IN2_i <= "00110100110010111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011101110";
   IN2_i <= "00110100111101101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101001100";
   IN2_i <= "00100101000011001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100100000";
   IN2_i <= "01000011011110010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100111101";
   IN2_i <= "00000000001010000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001011010";
   IN2_i <= "00001100000111001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111010110";
   IN2_i <= "00111010100010011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011000111";
   IN2_i <= "01111010011100100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010101011";
   IN2_i <= "00000110101000100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111011";
   IN2_i <= "00100010010100010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101100101";
   IN2_i <= "00111001011010111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010000010";
   IN2_i <= "00001110110101110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001101110";
   IN2_i <= "00011100001110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111001001";
   IN2_i <= "00010001001001011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101011111";
   IN2_i <= "00101101000001011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010110";
   IN2_i <= "00111001111010111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110111001";
   IN2_i <= "00111010111111100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010000101";
   IN2_i <= "01110000010011110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111010111";
   IN2_i <= "01110111111110110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010011";
   IN2_i <= "00000011001010010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111010101";
   IN2_i <= "00100100111100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100111011";
   IN2_i <= "01111100100000000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100101011";
   IN2_i <= "00100001000001100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101111001";
   IN2_i <= "01111111000011111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111110100";
   IN2_i <= "01110101011110011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011001011";
   IN2_i <= "01110010110100010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101011110";
   IN2_i <= "00010000001010000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111010010";
   IN2_i <= "00001110001101101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100100";
   IN2_i <= "00010010111000100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101110101";
   IN2_i <= "01101100001001001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111101101";
   IN2_i <= "01101011001000000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000110001";
   IN2_i <= "00110100001011010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000000101";
   IN2_i <= "01001110101001100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001111010";
   IN2_i <= "00011101010011100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001011000";
   IN2_i <= "01101101010010110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110110010";
   IN2_i <= "00001100110001001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101011111";
   IN2_i <= "00001111001101110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001010001";
   IN2_i <= "00010010101111111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010111000";
   IN2_i <= "01001000010000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000001010";
   IN2_i <= "00100110111010110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010001100";
   IN2_i <= "01011100101001011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110100100";
   IN2_i <= "00010000011101111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101101101";
   IN2_i <= "00010010100110011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100110010";
   IN2_i <= "00010110110100010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011111110";
   IN2_i <= "00101110111001000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011101001";
   IN2_i <= "00100101110010100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110101";
   IN2_i <= "00011011110010011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101010000";
   IN2_i <= "01111111011011110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100110101";
   IN2_i <= "01110110100101000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100111100";
   IN2_i <= "01010011011101110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101100011";
   IN2_i <= "00110001010000100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101000001";
   IN2_i <= "00110001001010110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001011100";
   IN2_i <= "01001101100011101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100001101";
   IN2_i <= "01111001111100000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101010";
   IN2_i <= "00011011011111000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011110000";
   IN2_i <= "01111110101000110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100110000";
   IN2_i <= "01011000001001100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001100101";
   IN2_i <= "01000110110011011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111111010";
   IN2_i <= "00110111101010010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000010100";
   IN2_i <= "00100101101100011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101000010";
   IN2_i <= "01111011101011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111001";
   IN2_i <= "01011011010111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000011100";
   IN2_i <= "00101000110011111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010011000";
   IN2_i <= "01101001010110011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100010001";
   IN2_i <= "00000100111101111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000011010";
   IN2_i <= "00110010111001001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011100101";
   IN2_i <= "00110100010010001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110000101";
   IN2_i <= "00000011011101001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000101011";
   IN2_i <= "00011011000001110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100101000";
   IN2_i <= "01001111110001011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011010";
   IN2_i <= "00010011000010100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110100101";
   IN2_i <= "00011010001011001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100110001";
   IN2_i <= "00000100010110110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100100001";
   IN2_i <= "00100000100001110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101011111";
   IN2_i <= "00110101100010101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100001";
   IN2_i <= "00111101101001001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011001111";
   IN2_i <= "01111010110011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111010010";
   IN2_i <= "01110100001011111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110000100";
   IN2_i <= "01110001111110111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100101110";
   IN2_i <= "00101101101111101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100111000";
   IN2_i <= "01111011011101101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001101010";
   IN2_i <= "00111110100001001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100011010";
   IN2_i <= "00010001111011000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011111110";
   IN2_i <= "01001101010111110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100000110";
   IN2_i <= "00100101010011100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110011011";
   IN2_i <= "00000000110101001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011100001";
   IN2_i <= "01011111011000100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011110101";
   IN2_i <= "00100000010101100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011111000";
   IN2_i <= "01100000110100111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100101111";
   IN2_i <= "00010111001001011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111010000";
   IN2_i <= "00111101111000111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010010000";
   IN2_i <= "01110010001111101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110010101";
   IN2_i <= "01001110001011111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011011111";
   IN2_i <= "00011110011000011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101001001";
   IN2_i <= "01110001100011110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000101101";
   IN2_i <= "01010110010010100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010011101";
   IN2_i <= "00001011101101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101110100";
   IN2_i <= "00010010001001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100110010";
   IN2_i <= "01001100111000100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111101000";
   IN2_i <= "00100111010001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001101111";
   IN2_i <= "00100011110010010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000111001";
   IN2_i <= "00011011111000110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010011111";
   IN2_i <= "01010101011101010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100010101";
   IN2_i <= "00111010110001001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100011100";
   IN2_i <= "00100011000111111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010110100";
   IN2_i <= "00000001000010011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011111000";
   IN2_i <= "00000000011110110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100011100";
   IN2_i <= "00001010011100001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001111";
   IN2_i <= "01110110011111000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100001000";
   IN2_i <= "00010000101010101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011100000";
   IN2_i <= "01100101010001010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111010011";
   IN2_i <= "01100111010101010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001111100";
   IN2_i <= "00011001111110000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001001101";
   IN2_i <= "00111001101000011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100010110";
   IN2_i <= "01100111111000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100000";
   IN2_i <= "00010011100110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100111101";
   IN2_i <= "01000110001010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010101001";
   IN2_i <= "01010111110111001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111000100";
   IN2_i <= "01000110010101100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000101011";
   IN2_i <= "00011101111001010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001101010";
   IN2_i <= "01001110011001110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001000001";
   IN2_i <= "01001001001000010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110000010";
   IN2_i <= "01010111100101001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101000011";
   IN2_i <= "00110000001101101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111111100";
   IN2_i <= "01000101111101011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100101111";
   IN2_i <= "00110100100011011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011010010";
   IN2_i <= "00111000001011100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001011101";
   IN2_i <= "00000101000101011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100110110";
   IN2_i <= "01011101000011011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100011001";
   IN2_i <= "01100011000100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110100001";
   IN2_i <= "00000100011100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100100100";
   IN2_i <= "01000110100001010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011111100";
   IN2_i <= "00011100101011001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101001011";
   IN2_i <= "00101111110101001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101101110";
   IN2_i <= "01011100111111001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110110000";
   IN2_i <= "01011100100001010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100110111";
   IN2_i <= "00100101011100111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101000101";
   IN2_i <= "00001000101011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101111000";
   IN2_i <= "01110111011100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010111110";
   IN2_i <= "00111000100001001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101100011";
   IN2_i <= "01001101001011100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001010011";
   IN2_i <= "00110001000001100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111000011";
   IN2_i <= "00111100110010011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100110100";
   IN2_i <= "01111111001000000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110110110";
   IN2_i <= "00011001011011011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111110000";
   IN2_i <= "00000110110000010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110111101";
   IN2_i <= "00110101101111101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111110010";
   IN2_i <= "01011101010011001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110011011";
   IN2_i <= "01000100001110000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111010110";
   IN2_i <= "00000011101100101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011111110";
   IN2_i <= "01111101111001101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110111101";
   IN2_i <= "01010011110100001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010011011";
   IN2_i <= "00101011111101110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100101010";
   IN2_i <= "01110000101110100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000111110";
   IN2_i <= "00101001110100101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001111101";
   IN2_i <= "00010000001000111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000000011";
   IN2_i <= "00100100001000010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011110001";
   IN2_i <= "01101001001111100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010011100";
   IN2_i <= "01110110011100011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011100";
   IN2_i <= "01110100100100100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110011000";
   IN2_i <= "01101011011011011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111100011";
   IN2_i <= "00011001111001100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111001111";
   IN2_i <= "00010111110001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001010010";
   IN2_i <= "01010011110110110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101010011";
   IN2_i <= "00010100010000010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011101101";
   IN2_i <= "01000101001001001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100010100";
   IN2_i <= "01111010000001010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000010101";
   IN2_i <= "00100100010001010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000110001";
   IN2_i <= "01101111000100010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111010011";
   IN2_i <= "01110111000011100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001010100";
   IN2_i <= "01001101110000111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010010011";
   IN2_i <= "01001101001000010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101000011";
   IN2_i <= "00100100100000010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001000111";
   IN2_i <= "01101001000000000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010000010";
   IN2_i <= "00000000110100011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111000010";
   IN2_i <= "01001101010011000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010001100";
   IN2_i <= "00001010011100100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001100001";
   IN2_i <= "00100111011000000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000111001";
   IN2_i <= "00011100110111101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010001011";
   IN2_i <= "01101000000010010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101000010";
   IN2_i <= "00101100001010000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100110";
   IN2_i <= "01000110100100101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011101000";
   IN2_i <= "01111011101010111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000100111";
   IN2_i <= "01000101011110010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011011000";
   IN2_i <= "00011011111011100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101000011";
   IN2_i <= "01000101011000010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101011011";
   IN2_i <= "01010011001111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111111011";
   IN2_i <= "00100011100101000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111010110";
   IN2_i <= "01001001110110111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111010111";
   IN2_i <= "00111010001100010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101010010";
   IN2_i <= "01101001001011100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011010011";
   IN2_i <= "01001100110010011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010001111";
   IN2_i <= "00100000001001101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111101001";
   IN2_i <= "01010110100010110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100011000";
   IN2_i <= "00010111010100110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110010111";
   IN2_i <= "01101110010111101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110000110";
   IN2_i <= "01011000010100101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011011101";
   IN2_i <= "00110000001101010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000000101";
   IN2_i <= "01010011100001111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000101011";
   IN2_i <= "00110010011000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101101011";
   IN2_i <= "01110011110111100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101001111";
   IN2_i <= "01001100010101011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101100001";
   IN2_i <= "00010111010000010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010110011";
   IN2_i <= "01111001101010111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101011111";
   IN2_i <= "00101100110100010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010010011";
   IN2_i <= "01001110001111111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111000101";
   IN2_i <= "01101001011010010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011101100";
   IN2_i <= "01110011110011000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111100100";
   IN2_i <= "00100101111101110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101110110";
   IN2_i <= "01001001000000001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101111001";
   IN2_i <= "01000001000011010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100010101";
   IN2_i <= "00001000000001111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100111010";
   IN2_i <= "00011011000011001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010010000";
   IN2_i <= "00000100011101111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000010010";
   IN2_i <= "00000000001100011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111101001";
   IN2_i <= "00010100110101110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010001";
   IN2_i <= "01101010001110011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000101110";
   IN2_i <= "01010100100011000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110000011";
   IN2_i <= "00000101011000101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101001011";
   IN2_i <= "01101101100010000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011000100";
   IN2_i <= "00000110001101011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111001010";
   IN2_i <= "00100100011111110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101101";
   IN2_i <= "01011011100111110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111001";
   IN2_i <= "00010011000111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010100001";
   IN2_i <= "00000001000010000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001110110";
   IN2_i <= "00111101100001001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000110010";
   IN2_i <= "00101100000011100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101010011";
   IN2_i <= "00101100011110111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110011011";
   IN2_i <= "00111000100111111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101010";
   IN2_i <= "00100010100001111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111001100";
   IN2_i <= "00100110010110001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011101010";
   IN2_i <= "00000101010110100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011010110";
   IN2_i <= "01010000110100101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101011001";
   IN2_i <= "00011111011100001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111001011";
   IN2_i <= "00001100101000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011000011";
   IN2_i <= "01001000101001101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011100001";
   IN2_i <= "01000101100011001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110110";
   IN2_i <= "00011111111000110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101110101";
   IN2_i <= "01010101110111011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101101000";
   IN2_i <= "00110101101111100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110010011";
   IN2_i <= "00101010000110111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100000110";
   IN2_i <= "01110010111000010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010101110";
   IN2_i <= "01111010000011100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110111101";
   IN2_i <= "00101010111000010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100011010";
   IN2_i <= "00000000001010011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000010010";
   IN2_i <= "00110100000100001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110101010";
   IN2_i <= "01011110011110110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011111011";
   IN2_i <= "00111111000110010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101101000";
   IN2_i <= "00000001100011010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101010";
   IN2_i <= "01001100001010010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011011110";
   IN2_i <= "00011011100101100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101111010";
   IN2_i <= "00100101011010011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110011101";
   IN2_i <= "00100000101010111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010100111";
   IN2_i <= "00010011100101000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011010011";
   IN2_i <= "00010100010000000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011110110";
   IN2_i <= "01110111011101100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110101";
   IN2_i <= "01100010101010111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010110010";
   IN2_i <= "01111001101000011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010001011";
   IN2_i <= "00101101110111101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001000010";
   IN2_i <= "00100010010010111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001100111";
   IN2_i <= "01000100110111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010000";
   IN2_i <= "00111100101010011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001111110";
   IN2_i <= "01011110111101010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111110100";
   IN2_i <= "00100011101111101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100000100";
   IN2_i <= "00011001000000101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010101";
   IN2_i <= "00111100000101110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110011110";
   IN2_i <= "01000001001101101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111000011";
   IN2_i <= "01110111011101101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010010010";
   IN2_i <= "00001101000110110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111001011";
   IN2_i <= "01110100101100100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001010111";
   IN2_i <= "00010011111000010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101101000";
   IN2_i <= "00111111101011110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001011111";
   IN2_i <= "00010000010001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100010000";
   IN2_i <= "00011100101101110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010000111";
   IN2_i <= "01111001110100000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010010";
   IN2_i <= "01001111001111010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100011";
   IN2_i <= "00010110110001101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101110011";
   IN2_i <= "00010000001001100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101010011";
   IN2_i <= "00010111011001110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110100110";
   IN2_i <= "01111101000101100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011110";
   IN2_i <= "00011011001011100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100100110";
   IN2_i <= "01111000110001111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101101";
   IN2_i <= "01000101110100011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100101001";
   IN2_i <= "00011111100011110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001111001";
   IN2_i <= "01001111101011111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000100011";
   IN2_i <= "00011100100010010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010001011";
   IN2_i <= "00001110111000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100010001";
   IN2_i <= "00011110101110100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100110100";
   IN2_i <= "00111100100111101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001010011";
   IN2_i <= "00100111110101010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001111010";
   IN2_i <= "01000000001111101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011111111";
   IN2_i <= "00111110101100011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000111110";
   IN2_i <= "01011111001101010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100110001";
   IN2_i <= "01100011100111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101101010";
   IN2_i <= "00011110011001011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011110010";
   IN2_i <= "01110110100011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011000110";
   IN2_i <= "00011110000110101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011100100";
   IN2_i <= "00000011110001000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001110010";
   IN2_i <= "01001011011010111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001001001";
   IN2_i <= "01110010011101101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011100";
   IN2_i <= "00010000011111110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010110100";
   IN2_i <= "00100000100010100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110010011";
   IN2_i <= "01011000100111001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010111111";
   IN2_i <= "01101000111010100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011000111";
   IN2_i <= "01011111000000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110111001";
   IN2_i <= "01101111001001000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111101011";
   IN2_i <= "01011000001101101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001101";
   IN2_i <= "01011001000011100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111000";
   IN2_i <= "01000011110101000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000011";
   IN2_i <= "01000101001011110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010111111";
   IN2_i <= "00000001111001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100110111";
   IN2_i <= "00000001100101011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110110";
   IN2_i <= "01110011101011010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111100110";
   IN2_i <= "00100011110111100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110010110";
   IN2_i <= "01101001100001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101110011";
   IN2_i <= "00110101101111100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110000010";
   IN2_i <= "01000011111000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011110111";
   IN2_i <= "00011110000011110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100101101";
   IN2_i <= "01011110100100000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111111111";
   IN2_i <= "00101101000001100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011001010";
   IN2_i <= "01111010101101001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111011";
   IN2_i <= "00101100111000110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001000";
   IN2_i <= "01001100001111110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010101011";
   IN2_i <= "00000001001000011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110011001";
   IN2_i <= "00111001011100011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000010010";
   IN2_i <= "00100111101111011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001000101";
   IN2_i <= "01101010100100110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111111101";
   IN2_i <= "00100011110000100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010111000";
   IN2_i <= "01000111110000000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101100001";
   IN2_i <= "00101110010001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110101";
   IN2_i <= "01101000010110111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001101000";
   IN2_i <= "01001001001011111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011001000";
   IN2_i <= "00010110011111011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100001111";
   IN2_i <= "01000101001010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111101110";
   IN2_i <= "00100100010110000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101001";
   IN2_i <= "00010010010010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100101010";
   IN2_i <= "01000000010000101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011100001";
   IN2_i <= "00101010101100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101111100";
   IN2_i <= "01100010111000101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011110010";
   IN2_i <= "01000101101010111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110011100";
   IN2_i <= "00101001000000100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110010101";
   IN2_i <= "00011100110011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100110111";
   IN2_i <= "01100100010010011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111001101";
   IN2_i <= "00011100001001110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101000010";
   IN2_i <= "01000000101000001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010111110";
   IN2_i <= "00100110000010000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111110101";
   IN2_i <= "00110111101110011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011001000";
   IN2_i <= "01011110010101010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110011010";
   IN2_i <= "01001111100111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001010110";
   IN2_i <= "01011001111110100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111011001";
   IN2_i <= "00010001001010001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011101110";
   IN2_i <= "01001111111110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100111100";
   IN2_i <= "00001001100000011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011011000";
   IN2_i <= "00100011010110100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100000110";
   IN2_i <= "01010101101010100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000110";
   IN2_i <= "01111110111000011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011000";
   IN2_i <= "00010011011110110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011011111";
   IN2_i <= "01010101010011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001000110";
   IN2_i <= "00111101001111011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000010100";
   IN2_i <= "00000001010000000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011000100";
   IN2_i <= "01000010000010110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011010001";
   IN2_i <= "00110100010100101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011001111";
   IN2_i <= "00000110000010101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100001";
   IN2_i <= "01000111100111100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000000001";
   IN2_i <= "00111101010101010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100011111";
   IN2_i <= "01100111011111001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110101101";
   IN2_i <= "01111000111110000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011111101";
   IN2_i <= "01010010000100111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110110010";
   IN2_i <= "00000010111010100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001001001";
   IN2_i <= "00001100111100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001101001";
   IN2_i <= "01011110001101111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000010000";
   IN2_i <= "00011010000001000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011100011";
   IN2_i <= "00100001010101111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000010000";
   IN2_i <= "01010000011010001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101010001";
   IN2_i <= "00010100001100010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100101001";
   IN2_i <= "00000010111010111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000010";
   IN2_i <= "01101010010100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011011010";
   IN2_i <= "00111110010000101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011010000";
   IN2_i <= "01011000111101000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011010011";
   IN2_i <= "01110110100111101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000011001";
   IN2_i <= "00000101111110110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100101001";
   IN2_i <= "01001001011010101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100000";
   IN2_i <= "00101000110110100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001000100";
   IN2_i <= "01011001101011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111110101";
   IN2_i <= "00110010011100110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011000110";
   IN2_i <= "00000110101101000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011000101";
   IN2_i <= "01001111011100101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010011111";
   IN2_i <= "00101000001010000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010011010";
   IN2_i <= "01010001011011011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110111";
   IN2_i <= "00110000111001000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100011111";
   IN2_i <= "01001110111100011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010000101";
   IN2_i <= "00010101010010000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011010111";
   IN2_i <= "01001110001011111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101110101";
   IN2_i <= "01000111011101000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001011101";
   IN2_i <= "00101000110101011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000100110";
   IN2_i <= "00111110011000101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000110111";
   IN2_i <= "01011110110011011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110010011";
   IN2_i <= "00101011101001001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000100010";
   IN2_i <= "01100101000110011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110010100";
   IN2_i <= "01011010010001111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000011010";
   IN2_i <= "01111111001111011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110000101";
   IN2_i <= "01110100010001101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101101001";
   IN2_i <= "00010011000110011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110001101";
   IN2_i <= "00101011100000111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010111100";
   IN2_i <= "01100110010100101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000110011";
   IN2_i <= "00000001010101111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000000110";
   IN2_i <= "00101111110101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010000100";
   IN2_i <= "00010110010010011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011000100";
   IN2_i <= "00011111011011101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001100011";
   IN2_i <= "00111111010111110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101011010";
   IN2_i <= "00100011011111111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100011111";
   IN2_i <= "01001101110100001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000111000";
   IN2_i <= "00101111101011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010101011";
   IN2_i <= "01110111001110111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011010";
   IN2_i <= "00011011101101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000011011";
   IN2_i <= "00110100011010000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100100011";
   IN2_i <= "01011011011011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111111101";
   IN2_i <= "01001101111010001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110010010";
   IN2_i <= "00110110110000000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010110101";
   IN2_i <= "00011101110111010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011110000";
   IN2_i <= "01100110100010101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010000010";
   IN2_i <= "01100100100001010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001101010";
   IN2_i <= "01010010111010010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111010110";
   IN2_i <= "00011001011111111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011001111";
   IN2_i <= "00011100010000000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001100000";
   IN2_i <= "01101110100110111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010101011";
   IN2_i <= "00111111101100010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101110000";
   IN2_i <= "01100101100110010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011100101";
   IN2_i <= "00101001101101100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101101000";
   IN2_i <= "00111100010100000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011111001";
   IN2_i <= "01111010001001010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011000001";
   IN2_i <= "00000110100000101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011011111";
   IN2_i <= "01001000011110000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001001";
   IN2_i <= "00000010111100011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110000111";
   IN2_i <= "01101001010110110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101001010";
   IN2_i <= "00010100011011001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001001111";
   IN2_i <= "00101111011000000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110011100";
   IN2_i <= "01111010100000000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010010101";
   IN2_i <= "00010010000001100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101110000";
   IN2_i <= "01011011001000000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110011011";
   IN2_i <= "01011101001010100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011000011";
   IN2_i <= "00010111100011000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010101000";
   IN2_i <= "00101110100010001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100101011";
   IN2_i <= "01001100111101110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110001101";
   IN2_i <= "01001111100011101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000001101";
   IN2_i <= "00000110100101011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111000010";
   IN2_i <= "01111011100010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011100100";
   IN2_i <= "01110011110101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000111111";
   IN2_i <= "01011001010010001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000001";
   IN2_i <= "01111000000100110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100111010";
   IN2_i <= "00110010000000111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010001101";
   IN2_i <= "00110010110010000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100011100";
   IN2_i <= "00000100101010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000011101";
   IN2_i <= "01101111101100010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101011001";
   IN2_i <= "00111001100111101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010101010";
   IN2_i <= "00011101010101111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010100100";
   IN2_i <= "01100110011110010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011110111";
   IN2_i <= "01010100111000111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101101110";
   IN2_i <= "01101010100001101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111010101";
   IN2_i <= "01101101101111101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110000";
   IN2_i <= "01001011000010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010100001";
   IN2_i <= "01101000001110110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111010110";
   IN2_i <= "01111001100001101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010100010";
   IN2_i <= "00010111011000000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011110101";
   IN2_i <= "00101111010110101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100110";
   IN2_i <= "01101100001011000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111111011";
   IN2_i <= "01100101011110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001010011";
   IN2_i <= "01000111110110100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110101";
   IN2_i <= "00110101111001100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001001101";
   IN2_i <= "01111010001111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100010110";
   IN2_i <= "00101000010110110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100101111";
   IN2_i <= "01100010111111011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101001011";
   IN2_i <= "00011101001111111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100001100";
   IN2_i <= "00000010101101000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011100110";
   IN2_i <= "00111110100100100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110111011";
   IN2_i <= "00100110010001100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000000010";
   IN2_i <= "01101111111010000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001001010";
   IN2_i <= "00011010110110101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100111111";
   IN2_i <= "01111110010110101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001010101";
   IN2_i <= "00100001000110010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101010001";
   IN2_i <= "00100001010010010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010111100";
   IN2_i <= "00110010111100000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101000010";
   IN2_i <= "01001000000111100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000011100";
   IN2_i <= "00101110111111001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000011010";
   IN2_i <= "01110100001100111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010010";
   IN2_i <= "01011100001111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011010111";
   IN2_i <= "00111001010111010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101110001";
   IN2_i <= "00011111001101110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101000010";
   IN2_i <= "01100110001110010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000111001";
   IN2_i <= "00100110100111100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111111";
   IN2_i <= "00101110101100010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100101100";
   IN2_i <= "01010011011101010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111111011";
   IN2_i <= "01101011100011110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110111010";
   IN2_i <= "00111100100110001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000011011";
   IN2_i <= "01101100100011000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111100111";
   IN2_i <= "00001100001101010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010101010";
   IN2_i <= "01011100111101010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111101111";
   IN2_i <= "01010001000010011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011010010";
   IN2_i <= "00111001000010000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110000111";
   IN2_i <= "00000010101001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111101";
   IN2_i <= "01111000110001100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011110100";
   IN2_i <= "01111110000001001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011001010";
   IN2_i <= "00001011011101010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000101010";
   IN2_i <= "01101001010011100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100100001";
   IN2_i <= "01100001011100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101110101";
   IN2_i <= "01001100111001011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110001001";
   IN2_i <= "00100010011001100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011001000";
   IN2_i <= "01010101000101111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101001100";
   IN2_i <= "00101010011010100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011101101";
   IN2_i <= "01101010100111100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101001010";
   IN2_i <= "01110011111010011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111100111";
   IN2_i <= "00100011111110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001011";
   IN2_i <= "01011010100100111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101100111";
   IN2_i <= "01001000101100011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010001101";
   IN2_i <= "01101011000010000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101111000";
   IN2_i <= "01010110011010100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101010011";
   IN2_i <= "00100100011011100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000001101";
   IN2_i <= "01111000011010100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110010101";
   IN2_i <= "01001000011101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011010100";
   IN2_i <= "01100010111111000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000100000";
   IN2_i <= "01011010001010101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010111001";
   IN2_i <= "01010101101010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001101000";
   IN2_i <= "01000010000101001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100101111";
   IN2_i <= "00000011000111111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011011010";
   IN2_i <= "01010110101101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011011111";
   IN2_i <= "00110001100011000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100110011";
   IN2_i <= "01100001101100010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110100110";
   IN2_i <= "00010000101110011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101110110";
   IN2_i <= "01011010110110100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110110";
   IN2_i <= "01010010100100000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011101111";
   IN2_i <= "01100000101101001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001011001";
   IN2_i <= "00100100100111110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001011110";
   IN2_i <= "01000111000100000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011100000";
   IN2_i <= "01011110111011011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111010010";
   IN2_i <= "00100001000001110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100000001";
   IN2_i <= "00111110011001100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000111000";
   IN2_i <= "00101011111111011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110011100";
   IN2_i <= "00110110000110001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010110011";
   IN2_i <= "00001110111101010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010110000";
   IN2_i <= "00111011011011010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111101110";
   IN2_i <= "01010101110101010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000010010";
   IN2_i <= "00101111101111111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110010000";
   IN2_i <= "00001010111100000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101000000";
   IN2_i <= "00010000011101001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001010";
   IN2_i <= "00100001110000011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010100100";
   IN2_i <= "00000111000011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000111000";
   IN2_i <= "00100101101111001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010111011";
   IN2_i <= "01111111100011011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110001101";
   IN2_i <= "00100110101110100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001101011";
   IN2_i <= "00001011111011100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011000010";
   IN2_i <= "01010010010001001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010100010";
   IN2_i <= "01100010000010011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101100";
   IN2_i <= "00110101011000100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100011110";
   IN2_i <= "00101010000011101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110101110";
   IN2_i <= "01111011001010000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101011010";
   IN2_i <= "01010111001011111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111010010";
   IN2_i <= "00001111111011101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011001110";
   IN2_i <= "01001010111110110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001110011";
   IN2_i <= "01011011111011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011111111";
   IN2_i <= "00000010111011100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110101111";
   IN2_i <= "01100101001011101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011010000";
   IN2_i <= "01001110111111111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110100010";
   IN2_i <= "01111001011101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011110111";
   IN2_i <= "00011000001110001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100101001";
   IN2_i <= "00101111010011101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111010000";
   IN2_i <= "00111111001110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101111100";
   IN2_i <= "01111101001101101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010000001";
   IN2_i <= "01000100001111000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011111000";
   IN2_i <= "00001111011111101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100000100";
   IN2_i <= "00001101001001110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000100000";
   IN2_i <= "01011010001110110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101000010";
   IN2_i <= "00010111010110101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110010100";
   IN2_i <= "01010011100011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001110010";
   IN2_i <= "01010101111000100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100110100";
   IN2_i <= "00000011001101001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101101001";
   IN2_i <= "00000111011000100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100001000";
   IN2_i <= "01000001001001100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101001111";
   IN2_i <= "00000011101100111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101011110";
   IN2_i <= "00110001001010111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100011110";
   IN2_i <= "00010010010110011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001100";
   IN2_i <= "00101110111011011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111011000";
   IN2_i <= "00110001001010010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101000001";
   IN2_i <= "01000101101011111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011101011";
   IN2_i <= "01000111110001111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011011000";
   IN2_i <= "00001111010001110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100110100";
   IN2_i <= "00001110111110000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000010010";
   IN2_i <= "01001101001011100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110110000";
   IN2_i <= "00000110110001110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000110101";
   IN2_i <= "00011001111010001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011100011";
   IN2_i <= "01101111100100001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010000101";
   IN2_i <= "01000000000000011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000000001";
   IN2_i <= "00000011001001101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101001001";
   IN2_i <= "01011001111110101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110111101";
   IN2_i <= "01010001100001101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010100000";
   IN2_i <= "01100001001111010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100010111";
   IN2_i <= "01110110100001100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111011011";
   IN2_i <= "01010100000000111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011011101";
   IN2_i <= "01111110000011101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010000011";
   IN2_i <= "00011110101111111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010011101";
   IN2_i <= "01100010001111111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101000110";
   IN2_i <= "01111101101010010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001001010";
   IN2_i <= "01101101110100011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101001011";
   IN2_i <= "01110011001111110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010011001";
   IN2_i <= "01110000101010100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101000101";
   IN2_i <= "01000100000111000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001111110";
   IN2_i <= "00000111110100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011001000";
   IN2_i <= "01001011011010111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001001011";
   IN2_i <= "01000011110110001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110111111";
   IN2_i <= "01010001011111101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101001110";
   IN2_i <= "01110011010110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100100000";
   IN2_i <= "00011111100010000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100011011";
   IN2_i <= "00011000001000111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011000011";
   IN2_i <= "00100100101101010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000110101";
   IN2_i <= "01100000100000111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111010001";
   IN2_i <= "01001010111000010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010111001";
   IN2_i <= "01110000011101010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010011110";
   IN2_i <= "00010000010000011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011000011";
   IN2_i <= "00000100010010111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000000101";
   IN2_i <= "01000110010010010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010110000";
   IN2_i <= "01010111010100010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010011010";
   IN2_i <= "01000101011110011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100011010";
   IN2_i <= "00100001101110010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101000100";
   IN2_i <= "00011011110111101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000100001";
   IN2_i <= "00110111000000101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110100";
   IN2_i <= "00001000010010001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010000110";
   IN2_i <= "00101000100110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001011101";
   IN2_i <= "01010111000100000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001001101";
   IN2_i <= "00101011011001011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111110011";
   IN2_i <= "01100000000001000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111100010";
   IN2_i <= "00110010100111001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010010101";
   IN2_i <= "01010101100010101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111001000";
   IN2_i <= "00111011010100000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101110";
   IN2_i <= "00100001111010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000110011";
   IN2_i <= "01110101000100101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101000010";
   IN2_i <= "00010111101011101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100101100";
   IN2_i <= "00100100100011000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001010000";
   IN2_i <= "00010100110000101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011010000";
   IN2_i <= "01010111011111000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010011010";
   IN2_i <= "00100000011111110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010110010";
   IN2_i <= "01110010110011010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111010101";
   IN2_i <= "01110100100001001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111000011";
   IN2_i <= "00000001011111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101010011";
   IN2_i <= "00110100111011001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000111100";
   IN2_i <= "00010011000010101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100010100";
   IN2_i <= "01100000110000010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100101100";
   IN2_i <= "01000000001100100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010011100";
   IN2_i <= "01100101001100100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110010110";
   IN2_i <= "01001011110100001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110010111";
   IN2_i <= "00111001100101101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010011011";
   IN2_i <= "00100010110110000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011001";
   IN2_i <= "01010011010000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111001010";
   IN2_i <= "00000000110011001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010101001";
   IN2_i <= "01000011100110101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110000111";
   IN2_i <= "00000010110101001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100110111";
   IN2_i <= "01010100000000110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100010011";
   IN2_i <= "00000010100010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110110001";
   IN2_i <= "01101111010110100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100111011";
   IN2_i <= "00101000101011101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001011";
   IN2_i <= "00100001111111000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010101";
   IN2_i <= "01110101100010111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011100001";
   IN2_i <= "00010111111111111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101111";
   IN2_i <= "01100110111000101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000011";
   IN2_i <= "00100001111111001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000010110";
   IN2_i <= "01011101001100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101000010";
   IN2_i <= "01110011111000100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110111110";
   IN2_i <= "00001000100100100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101110";
   IN2_i <= "00011000001010001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000101010";
   IN2_i <= "00010011100110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011001000";
   IN2_i <= "00000010111111011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000010111";
   IN2_i <= "01100010011101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100100000";
   IN2_i <= "01011111100100010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100110100";
   IN2_i <= "00011111100000011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110010011";
   IN2_i <= "00011010000011110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011101110";
   IN2_i <= "00111101011011011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010000000";
   IN2_i <= "00010001110000010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000100000";
   IN2_i <= "01000110001000011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111110110";
   IN2_i <= "00011101010110111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010110100";
   IN2_i <= "01011011111101100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001100000";
   IN2_i <= "01100011111010011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101100101";
   IN2_i <= "01000000100011000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100100001";
   IN2_i <= "00001000010110101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110101100";
   IN2_i <= "01001000111101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011010111";
   IN2_i <= "01010101100100011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111010110";
   IN2_i <= "01110011100100011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111001";
   IN2_i <= "00101111010010111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100110110";
   IN2_i <= "00110110000100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011100010";
   IN2_i <= "00110001010010011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001001111";
   IN2_i <= "01010101111100001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011011100";
   IN2_i <= "01000001110011111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010011011";
   IN2_i <= "00100101101000001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000111101";
   IN2_i <= "00101111111001011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100000111";
   IN2_i <= "01100111101000000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100011010";
   IN2_i <= "00100011111000100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001001000";
   IN2_i <= "01110001111110101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001011101";
   IN2_i <= "01101110110101100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000011100";
   IN2_i <= "00100010111001010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111010000";
   IN2_i <= "00110100111101010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100100";
   IN2_i <= "01110111110011001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010110";
   IN2_i <= "01110100001011100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000010100";
   IN2_i <= "01101010010111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010001101";
   IN2_i <= "00011111000111100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101101000";
   IN2_i <= "01011000110010010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101001000";
   IN2_i <= "01101011101010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100000110";
   IN2_i <= "00001100110101100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001011011";
   IN2_i <= "01011011011110111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101110011";
   IN2_i <= "00110011101011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101010100";
   IN2_i <= "01110000101011000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010001011";
   IN2_i <= "00011010011110010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010111010";
   IN2_i <= "01111101000011100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000000010";
   IN2_i <= "00011101111111010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111000011";
   IN2_i <= "01111101010001100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111001011";
   IN2_i <= "01111110101010111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010000100";
   IN2_i <= "01010100110110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110110011";
   IN2_i <= "01101110100011011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101011111";
   IN2_i <= "00100011100100111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100110100";
   IN2_i <= "00101000000111001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010110101";
   IN2_i <= "00101101100100010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011100100";
   IN2_i <= "01101000001101111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110000000";
   IN2_i <= "00111001000110100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101010110";
   IN2_i <= "00000100100100010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001010111";
   IN2_i <= "00011100101111111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100011100";
   IN2_i <= "01000000010100111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000001000";
   IN2_i <= "01101011001001100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011011110";
   IN2_i <= "00011000001000100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011010011";
   IN2_i <= "01110000010001000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010011010";
   IN2_i <= "00110001011010100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011010010";
   IN2_i <= "01011001111100101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100101000";
   IN2_i <= "00010101001000100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101110111";
   IN2_i <= "01100011010110001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110010100";
   IN2_i <= "01010011000111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010000010";
   IN2_i <= "00100110001111010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101011010";
   IN2_i <= "00011101101101101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100101000";
   IN2_i <= "01101011011111101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110011100";
   IN2_i <= "00000110110000111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100101011";
   IN2_i <= "00111010110110100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111011110";
   IN2_i <= "01101000000001100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001011110";
   IN2_i <= "01101100010100010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101000110";
   IN2_i <= "01000100111101010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001111010";
   IN2_i <= "01101010100110010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010010001";
   IN2_i <= "01110000000010100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110001000";
   IN2_i <= "01111001001011011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001111001";
   IN2_i <= "00111000110100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101001100";
   IN2_i <= "00011011111100100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011100000";
   IN2_i <= "01001101111100110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010010110";
   IN2_i <= "00101101110000000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110111100";
   IN2_i <= "01101110000111111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011011001";
   IN2_i <= "00101111101010110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001011100";
   IN2_i <= "00101001111000110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010101001";
   IN2_i <= "01010010010010111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100100010";
   IN2_i <= "01111110101100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100000110";
   IN2_i <= "01111111000111000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110101011";
   IN2_i <= "01100010100111010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001010011";
   IN2_i <= "00010111001010000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100111000";
   IN2_i <= "01001100111010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000000110";
   IN2_i <= "01000011011111001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100100000";
   IN2_i <= "00100111010101110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010111101";
   IN2_i <= "00000010111000101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100000110";
   IN2_i <= "00100011001010111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001001000";
   IN2_i <= "00100011111110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100000010";
   IN2_i <= "01101001110111101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000110001";
   IN2_i <= "01110000001110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000001010";
   IN2_i <= "01100100000011011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100100001";
   IN2_i <= "00010010010010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011101111";
   IN2_i <= "01000011001011100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011011100";
   IN2_i <= "00001101001101110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100101";
   IN2_i <= "00100000001111000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101011100";
   IN2_i <= "00011001101010101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000111111";
   IN2_i <= "01000001111000000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010110011";
   IN2_i <= "01001111001111011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101110";
   IN2_i <= "00010101010011010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011110001";
   IN2_i <= "01011010111010011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100101";
   IN2_i <= "01000111101101111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101100011";
   IN2_i <= "01010111100010100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101001101";
   IN2_i <= "01100010101100101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011000011";
   IN2_i <= "00101010011111101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111011110";
   IN2_i <= "00011001110001001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000110011";
   IN2_i <= "00001001111110101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110000001";
   IN2_i <= "01000110100101000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111110010";
   IN2_i <= "01001001110110111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011010000";
   IN2_i <= "01101000101111100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001010000";
   IN2_i <= "00100100110100011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101101000";
   IN2_i <= "01011100001011000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001001101";
   IN2_i <= "00100110010001110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000001110";
   IN2_i <= "01010010100111111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101000";
   IN2_i <= "01000001110011110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110010010";
   IN2_i <= "01111000100111111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110001001";
   IN2_i <= "01101110111110110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110100101";
   IN2_i <= "01001101110111111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100000001";
   IN2_i <= "01110001101110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000101011";
   IN2_i <= "00000110111010101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001011001";
   IN2_i <= "01000000100100110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000110000";
   IN2_i <= "01110111101010110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001011110";
   IN2_i <= "00101010000010111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111110001";
   IN2_i <= "01110001011101010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101011111";
   IN2_i <= "00001001101111000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011100011";
   IN2_i <= "00100100111001110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001111001";
   IN2_i <= "01100101011010000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011110101";
   IN2_i <= "00001110000000110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001111011";
   IN2_i <= "00011111001000010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010010001";
   IN2_i <= "00010000100001011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111100111";
   IN2_i <= "00000100101010011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101011";
   IN2_i <= "00001111011111001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011110001";
   IN2_i <= "00000100000100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110011101";
   IN2_i <= "00111110001110011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111010100";
   IN2_i <= "01000010111111101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001000111";
   IN2_i <= "01110000010101111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101001000";
   IN2_i <= "01000000000101111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010011011";
   IN2_i <= "01000001100100101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111000110";
   IN2_i <= "01110101001101110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101110011";
   IN2_i <= "00110110011110010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100001001";
   IN2_i <= "00010101010101111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101000100";
   IN2_i <= "01110001100000001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000110100";
   IN2_i <= "00111011100111110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110001001";
   IN2_i <= "00100111001001010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001111";
   IN2_i <= "01001111110110011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100111";
   IN2_i <= "01100111110101110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001101010";
   IN2_i <= "01101011010110001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110101011";
   IN2_i <= "01101000011100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000001101";
   IN2_i <= "01101010101000000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000001011";
   IN2_i <= "01110110000000001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011101010";
   IN2_i <= "00000101111101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011111010";
   IN2_i <= "00010000100011110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100110111";
   IN2_i <= "01001011001001111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101010111";
   IN2_i <= "00010000011000011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011010100";
   IN2_i <= "01101001010111011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100111";
   IN2_i <= "01100101111011100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101100";
   IN2_i <= "01010110010011000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010011010";
   IN2_i <= "01101010010011111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100110";
   IN2_i <= "01100100011111101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000011110";
   IN2_i <= "01011100011110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101100101";
   IN2_i <= "00000111001010101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010110000";
   IN2_i <= "01000010010000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001110111";
   IN2_i <= "01001001000010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011011101";
   IN2_i <= "01110000000011110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100011110";
   IN2_i <= "01100001000101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010101";
   IN2_i <= "01011000110101010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010000000";
   IN2_i <= "01000011011101110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110010011";
   IN2_i <= "01100100001000110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110011000";
   IN2_i <= "00111110001101110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011000100";
   IN2_i <= "00011011101101111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010101101";
   IN2_i <= "00001110111111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001101010";
   IN2_i <= "00111111011111001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011010111";
   IN2_i <= "00011110000000010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001011011";
   IN2_i <= "00011000010111110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111110100";
   IN2_i <= "01111001001010010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000100000";
   IN2_i <= "00100101000100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110011101";
   IN2_i <= "00001100001100010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110100110";
   IN2_i <= "00000010000100100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100010011";
   IN2_i <= "00011010111110001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010010110";
   IN2_i <= "00111011010100011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110001011";
   IN2_i <= "00110000010111001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101011000";
   IN2_i <= "01010011000000100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010110110";
   IN2_i <= "01110000001110100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100001";
   IN2_i <= "00011111011101111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101000110";
   IN2_i <= "01111011000011001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100011010";
   IN2_i <= "01000111001011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001110111";
   IN2_i <= "01001100001000011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010111101";
   IN2_i <= "01100111000101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110011011";
   IN2_i <= "00001100011011001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111101101";
   IN2_i <= "00101110001010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011011011";
   IN2_i <= "00001011111100111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010111";
   IN2_i <= "00001001011101100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001111010";
   IN2_i <= "01010111111010100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100100110";
   IN2_i <= "00000110010101101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101101100";
   IN2_i <= "00110100001001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011100011";
   IN2_i <= "00111001001100011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000010101";
   IN2_i <= "01000100111001011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001011000";
   IN2_i <= "01111000101101011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001010101";
   IN2_i <= "00011110100011110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010110001";
   IN2_i <= "01111111100001110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011100010";
   IN2_i <= "00110011000010100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101010111";
   IN2_i <= "00011001011100110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000101000";
   IN2_i <= "00000111001000101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111001100";
   IN2_i <= "00100111010010100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000110110";
   IN2_i <= "00101011110111000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110011010";
   IN2_i <= "01100110111100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010000100";
   IN2_i <= "00111111101110100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100110010";
   IN2_i <= "01100010000011001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000101100";
   IN2_i <= "00011110101011000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011001011";
   IN2_i <= "00011011011001110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001001010";
   IN2_i <= "00000001111110100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100011110";
   IN2_i <= "00010111100110001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110111111";
   IN2_i <= "00110000110011000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101101011";
   IN2_i <= "00000110010001011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011100010";
   IN2_i <= "00100011000101001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000011010";
   IN2_i <= "00100011011000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100111110";
   IN2_i <= "01011101001111001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110001111";
   IN2_i <= "01111110011111010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001110111";
   IN2_i <= "00010110101000110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100011110";
   IN2_i <= "00100001110101001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000111010";
   IN2_i <= "00101001000010010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010110101";
   IN2_i <= "00001001010011101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000000111";
   IN2_i <= "00011001000100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111001001";
   IN2_i <= "01110110111101001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101110101";
   IN2_i <= "01111000011101010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100001111";
   IN2_i <= "01001001111010011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101001";
   IN2_i <= "01101111101011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100011110";
   IN2_i <= "01101101111010010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101110000";
   IN2_i <= "01011110001100010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000011010";
   IN2_i <= "00011100000000101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101101011";
   IN2_i <= "00010100010011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010010110";
   IN2_i <= "00101011000110000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001111000";
   IN2_i <= "01000010011100101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010101110";
   IN2_i <= "00110011101010001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010001000";
   IN2_i <= "01111010011011100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011110101";
   IN2_i <= "00010110100110011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101110101";
   IN2_i <= "00010000010101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100110010";
   IN2_i <= "01100111010101001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110110000";
   IN2_i <= "00000100110110010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000111010";
   IN2_i <= "01101100010111100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000011110";
   IN2_i <= "00011100011000000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111101100";
   IN2_i <= "00101101000011110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001101101";
   IN2_i <= "01001101010100110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111111110";
   IN2_i <= "00100000000100000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001100101";
   IN2_i <= "00011010010100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101110011";
   IN2_i <= "00101100011010001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111101111";
   IN2_i <= "00000000110010100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100011011";
   IN2_i <= "00001010110110011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000111110";
   IN2_i <= "01011000110000100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001001000";
   IN2_i <= "00011010110010100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100110010";
   IN2_i <= "00000010010000110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100100111";
   IN2_i <= "00011011100001001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011000";
   IN2_i <= "00110100111010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101010010";
   IN2_i <= "00111011101011011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000111011";
   IN2_i <= "00110101110001110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001000000";
   IN2_i <= "01010001011011101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100001";
   IN2_i <= "01101101101110110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011110010";
   IN2_i <= "00110011001111010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011100101";
   IN2_i <= "00110010110110101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110010001";
   IN2_i <= "01111010110001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111100";
   IN2_i <= "00011101110000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001110010";
   IN2_i <= "00011010101000110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101000";
   IN2_i <= "00110110001101010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110110011";
   IN2_i <= "01001100100101001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000101111";
   IN2_i <= "00010011011111001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110001111";
   IN2_i <= "01010100010100000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001100110";
   IN2_i <= "00111100100010001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000101000";
   IN2_i <= "01010011000010001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001100110";
   IN2_i <= "01011000000001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000101100";
   IN2_i <= "00000011101101011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001101001";
   IN2_i <= "00011100100000111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000110110";
   IN2_i <= "01111100011011001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111001";
   IN2_i <= "00010110011010010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011000011";
   IN2_i <= "00101011100001100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000001011";
   IN2_i <= "01111111010110110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111010000";
   IN2_i <= "01000000001000111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010100110";
   IN2_i <= "01111100001101111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111111";
   IN2_i <= "00010010111001101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100100111";
   IN2_i <= "00011100110001011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010100101";
   IN2_i <= "01011101001000100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101110";
   IN2_i <= "01100110011001011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111101110";
   IN2_i <= "00110101111101111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011100111";
   IN2_i <= "01011001000000001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010011000";
   IN2_i <= "01000110100001000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100000011";
   IN2_i <= "00110100001010100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001110011";
   IN2_i <= "00110010001100101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000111001";
   IN2_i <= "00101110110111110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100011010";
   IN2_i <= "01111111101010010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000101110";
   IN2_i <= "00001000000100101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100110000";
   IN2_i <= "00001000000110011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110010101";
   IN2_i <= "01100000110000110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010100111";
   IN2_i <= "00000111111100100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000000100";
   IN2_i <= "00000011101110111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110110011";
   IN2_i <= "01101101111100101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110101110";
   IN2_i <= "00000010011101011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100101";
   IN2_i <= "01000010100010001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111101";
   IN2_i <= "01001111001011110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010110001";
   IN2_i <= "00101110011010100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011100111";
   IN2_i <= "00101101001111010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011110001";
   IN2_i <= "01101110010100001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000111101";
   IN2_i <= "01110100000100101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100111101";
   IN2_i <= "01100101011010001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111110";
   IN2_i <= "01001110001001010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110110";
   IN2_i <= "01101110100010001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101101000";
   IN2_i <= "01110011110110100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000110010";
   IN2_i <= "01011001100000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100101011";
   IN2_i <= "01111010001011001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010000101";
   IN2_i <= "01011110000011001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101001011";
   IN2_i <= "00010011111000001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110000011";
   IN2_i <= "01001001111110111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110100000";
   IN2_i <= "00000010111110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111010010";
   IN2_i <= "01010011000100110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000011000";
   IN2_i <= "01111111111111111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101101000";
   IN2_i <= "01111111101010000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001011100";
   IN2_i <= "00110110000110000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100000";
   IN2_i <= "01100110011010011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101001011";
   IN2_i <= "01000101101011000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001011000";
   IN2_i <= "01011110011101110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110111111";
   IN2_i <= "01011101010110110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110000";
   IN2_i <= "01011010100111000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010010";
   IN2_i <= "01000110101111100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011110111";
   IN2_i <= "01111111011010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000010111";
   IN2_i <= "01111100100111000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000011000";
   IN2_i <= "01011011001001111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111011010";
   IN2_i <= "00110100000110101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000001011";
   IN2_i <= "00111111110110011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000110011";
   IN2_i <= "00110011111110101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100011111";
   IN2_i <= "01001111111111000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010010010";
   IN2_i <= "01001001111111000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001111101";
   IN2_i <= "00011111111011010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011101001";
   IN2_i <= "01110100111111010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000000110";
   IN2_i <= "01011001110001000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001110110";
   IN2_i <= "00001000000000010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010000111";
   IN2_i <= "01111100001000000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110110010";
   IN2_i <= "00011011110101100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101001111";
   IN2_i <= "01001101001110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011110000";
   IN2_i <= "00100100100001001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011011101";
   IN2_i <= "00100111111001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010011100";
   IN2_i <= "00010100011001111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011101000";
   IN2_i <= "01110100110010010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010110011";
   IN2_i <= "00000101110101111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000101111";
   IN2_i <= "00010101001110000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011111010";
   IN2_i <= "01010011100100001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010111000";
   IN2_i <= "00001001001110010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111100";
   IN2_i <= "01011011010100110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110000010";
   IN2_i <= "01100000011110011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111110100";
   IN2_i <= "00101101001110101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001111011";
   IN2_i <= "00101011010111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101010011";
   IN2_i <= "01000000011011011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100000111";
   IN2_i <= "00001001101101100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101111100";
   IN2_i <= "00100101001001011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100100001";
   IN2_i <= "01100011000011010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111110001";
   IN2_i <= "01101001111111001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011100100";
   IN2_i <= "01010111110111100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100111001";
   IN2_i <= "01011011101011100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100111000";
   IN2_i <= "01010000000111101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001110001";
   IN2_i <= "00011101011001110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111001000";
   IN2_i <= "01101100101001111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111001011";
   IN2_i <= "00001011010100010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111111000";
   IN2_i <= "01111110000110011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000100010";
   IN2_i <= "00011100111010110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100000100";
   IN2_i <= "00110111100101000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100001010";
   IN2_i <= "00101100000000111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011111010";
   IN2_i <= "01101110111100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110111011";
   IN2_i <= "00011111101111000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000100000";
   IN2_i <= "01100100101010111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011111001";
   IN2_i <= "01010011000101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110011010";
   IN2_i <= "01101001001100101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111010010";
   IN2_i <= "01111000110111011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011011000";
   IN2_i <= "00111000001010110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111100000";
   IN2_i <= "00101000110000011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001010101";
   IN2_i <= "00000001100111010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110001101";
   IN2_i <= "00100000010110100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101011110";
   IN2_i <= "00011111110001000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101001110";
   IN2_i <= "00010011001111111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000010101";
   IN2_i <= "00000100111010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101011110";
   IN2_i <= "00101000010101101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000101";
   IN2_i <= "00111011011000110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010110100";
   IN2_i <= "00011111001110001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000011010";
   IN2_i <= "00110101111101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010000111";
   IN2_i <= "00110001001011111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001000110";
   IN2_i <= "01011011111011101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010100100";
   IN2_i <= "00000010010101110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100100010";
   IN2_i <= "00110100000011000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011000010";
   IN2_i <= "01001110101100110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001111010";
   IN2_i <= "00110111110010010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000011110";
   IN2_i <= "01000100011110110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110011111";
   IN2_i <= "00111010100000010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110010101";
   IN2_i <= "00111101010010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100110010";
   IN2_i <= "00010111101011001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100110101";
   IN2_i <= "01011001110100001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110011";
   IN2_i <= "01110100101111001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000000101";
   IN2_i <= "01111100001001100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100011000";
   IN2_i <= "01110111110011001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100001001";
   IN2_i <= "01011111111000110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000001010";
   IN2_i <= "01000101001010011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100010001";
   IN2_i <= "01110111111111111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000011011";
   IN2_i <= "00100011111010110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000010101";
   IN2_i <= "01111101001101110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011110000";
   IN2_i <= "00110100110000011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001101010";
   IN2_i <= "01011111010110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101101011";
   IN2_i <= "01101111111010011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011110000";
   IN2_i <= "00000110010100011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000111110";
   IN2_i <= "00110000110101000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011011011";
   IN2_i <= "00000101011000111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101110100";
   IN2_i <= "01011101000110001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001101010";
   IN2_i <= "01010001111101111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001101111";
   IN2_i <= "00001001111111011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000101000";
   IN2_i <= "00101010011101110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010011000";
   IN2_i <= "00011001000111110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011101100";
   IN2_i <= "01100110010111000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111010011";
   IN2_i <= "00010011100110101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011010000";
   IN2_i <= "00110110011000110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011000101";
   IN2_i <= "00001110111011011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010111001";
   IN2_i <= "01110101100010011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010110010";
   IN2_i <= "01000010100000001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001011110";
   IN2_i <= "00001011000001111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100100011";
   IN2_i <= "01110000010000010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010001";
   IN2_i <= "00010000111010101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001100100";
   IN2_i <= "00100011000111010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010110101";
   IN2_i <= "01100000010101001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011010000";
   IN2_i <= "00011101111010111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001110111";
   IN2_i <= "00101001001011000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011010100";
   IN2_i <= "01111100010011001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011111011";
   IN2_i <= "01010001000111101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000100110";
   IN2_i <= "01100001011010011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001010110";
   IN2_i <= "00011101001110010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111100001";
   IN2_i <= "01001100000001000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000011001";
   IN2_i <= "01111001000110101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111101110";
   IN2_i <= "00111011100100101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011001001";
   IN2_i <= "01101101000111100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000101110";
   IN2_i <= "00111101111011010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101100101";
   IN2_i <= "01001110011011101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110011001";
   IN2_i <= "00010010100101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001100010";
   IN2_i <= "00111010101000101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100000110";
   IN2_i <= "01111010100100100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010111101";
   IN2_i <= "01101010101001111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000110001";
   IN2_i <= "00111011011110111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100010001";
   IN2_i <= "00110000011011110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000001001";
   IN2_i <= "01110011001100100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111101";
   IN2_i <= "00100101001101101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011010100";
   IN2_i <= "00001010110100010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010110011";
   IN2_i <= "01011000111111101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011001000";
   IN2_i <= "01100101100111001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010111000";
   IN2_i <= "01010000000110101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101010010";
   IN2_i <= "00100000110000110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001101101";
   IN2_i <= "00101001010000001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011001011";
   IN2_i <= "00110001010111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110100000";
   IN2_i <= "01111111001011010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100100011";
   IN2_i <= "01001010011100011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111111111";
   IN2_i <= "01001110110000011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000110";
   IN2_i <= "01110011001011010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100110101";
   IN2_i <= "00000111100111111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111001101";
   IN2_i <= "00111100011101011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011000101";
   IN2_i <= "00100101110110000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101000111";
   IN2_i <= "01101001110000011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010101001";
   IN2_i <= "01010100000000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010100000";
   IN2_i <= "01001100101010100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011101101";
   IN2_i <= "00011011010011010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101111010";
   IN2_i <= "01010101110101001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010101110";
   IN2_i <= "00111011010011101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011000110";
   IN2_i <= "01101101101111100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001111111";
   IN2_i <= "01000101111000101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110111000";
   IN2_i <= "01111111001100100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001111111";
   IN2_i <= "01101111110110001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101000111";
   IN2_i <= "00011010001100110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111001100";
   IN2_i <= "00111000101011101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000010011";
   IN2_i <= "01111110000111110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101100000";
   IN2_i <= "01110001011001101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111101011";
   IN2_i <= "01010011101010000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010010101";
   IN2_i <= "00000000000101110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001000000";
   IN2_i <= "00011011000111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100111001";
   IN2_i <= "01010110111010100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010101111";
   IN2_i <= "01100010101011100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101110000";
   IN2_i <= "01001011110010111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011001111";
   IN2_i <= "01010100110000110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011110011";
   IN2_i <= "00011101010001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101010110";
   IN2_i <= "00110100110010100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001000100";
   IN2_i <= "01101100111100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001101111";
   IN2_i <= "01100010010100010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001101111";
   IN2_i <= "01000101100111111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000110101";
   IN2_i <= "00101000111111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000111010";
   IN2_i <= "00010100110000011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010100100";
   IN2_i <= "01101100111001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111101101";
   IN2_i <= "00101100111011011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100001010";
   IN2_i <= "01010111100011110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110000011";
   IN2_i <= "00110110000001000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011110111";
   IN2_i <= "01010110100100001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110111100";
   IN2_i <= "00100010010100001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000000";
   IN2_i <= "01101110110111001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110101001";
   IN2_i <= "00000001110010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100110000";
   IN2_i <= "00010011011100101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010011001";
   IN2_i <= "01110101110010101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110100111";
   IN2_i <= "01011110111011000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111111011";
   IN2_i <= "01011111010000110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010010010";
   IN2_i <= "00001111001000101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111001";
   IN2_i <= "01110011011000100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110010111";
   IN2_i <= "00010000110110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110110000";
   IN2_i <= "00111001000001100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000011101";
   IN2_i <= "00010011000110100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101000";
   IN2_i <= "00011001010111111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011001111";
   IN2_i <= "01010111011100010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010110010";
   IN2_i <= "00110100110011100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010110100";
   IN2_i <= "00011010010101001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001000001";
   IN2_i <= "01010010000101100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110111011";
   IN2_i <= "01001101110001100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001101001";
   IN2_i <= "01011010111101100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101100111";
   IN2_i <= "01100001001000101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011110110";
   IN2_i <= "00111110111101010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010010101";
   IN2_i <= "00111111000111001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100110010";
   IN2_i <= "00110001000111011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001010110";
   IN2_i <= "00101010110010101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011011000";
   IN2_i <= "00101000111111000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001111110";
   IN2_i <= "01110101110000101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011110011";
   IN2_i <= "00100101011110010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101100001";
   IN2_i <= "00111110101110010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000100010";
   IN2_i <= "01111000110100000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011111";
   IN2_i <= "00110000101101101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111000001";
   IN2_i <= "00010111011010011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110011100";
   IN2_i <= "00111101000111001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001110110";
   IN2_i <= "01110110000010011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101011000";
   IN2_i <= "01100000101110000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101001101";
   IN2_i <= "01100111100010111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011111111";
   IN2_i <= "00001011011000011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110111";
   IN2_i <= "00010111000100000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000101010";
   IN2_i <= "00110101100010111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100001111";
   IN2_i <= "01101100000011011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101110011";
   IN2_i <= "00011100011101110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011010";
   IN2_i <= "01101001010100011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111101010";
   IN2_i <= "00001010001001011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110011110";
   IN2_i <= "01011001101101011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111011";
   IN2_i <= "01100000100111111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010101100";
   IN2_i <= "01010001111100111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011111010";
   IN2_i <= "00011100110110110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111010110";
   IN2_i <= "00001111000000100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000111001";
   IN2_i <= "00001010100000101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100001010";
   IN2_i <= "01110011000110111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101001010";
   IN2_i <= "00111001111111100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011110001";
   IN2_i <= "00101111100100001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010011011";
   IN2_i <= "00111010000011110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100011000";
   IN2_i <= "00101110001110001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011010110";
   IN2_i <= "00100111010000001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011001011";
   IN2_i <= "00111001001110010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111100111";
   IN2_i <= "00010010010010010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110000";
   IN2_i <= "01000111101000100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111001101";
   IN2_i <= "00100011000110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000010011";
   IN2_i <= "01011101010011111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000100001";
   IN2_i <= "00000010010110010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001101000";
   IN2_i <= "00100110000110011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001000001";
   IN2_i <= "00101111101110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000101000";
   IN2_i <= "01101111100101111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000101100";
   IN2_i <= "01001110010101111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101010110";
   IN2_i <= "01011110111101110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011010110";
   IN2_i <= "01000100100000001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101001";
   IN2_i <= "01110000110010100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100001001";
   IN2_i <= "00110101001110010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010000";
   IN2_i <= "00110010100101011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100011001";
   IN2_i <= "00001111001110010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101011000";
   IN2_i <= "00100000110101010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010011100";
   IN2_i <= "01010101000101101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011000011";
   IN2_i <= "00101110100001001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111101000";
   IN2_i <= "01001001101011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001100010";
   IN2_i <= "01001010000110111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011101011";
   IN2_i <= "00101111100101111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100001";
   IN2_i <= "01101011101001001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000101011";
   IN2_i <= "00010110000111100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111110";
   IN2_i <= "01000011110000110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100110111";
   IN2_i <= "00101001011000111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111111101";
   IN2_i <= "00100100110011111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100011001";
   IN2_i <= "01100100001010010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111001";
   IN2_i <= "01100011011101101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001110010";
   IN2_i <= "01010010110110111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010111010";
   IN2_i <= "01101000101110110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000001110";
   IN2_i <= "00110111101011010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000101110";
   IN2_i <= "00100011010001111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010100011";
   IN2_i <= "01101010100101000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111110111";
   IN2_i <= "01100010011110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011100110";
   IN2_i <= "01100101100010001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011011110";
   IN2_i <= "01000100101011110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000100011";
   IN2_i <= "00110001100101011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100011010";
   IN2_i <= "01010001000001010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010100011";
   IN2_i <= "00100001110000110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000110100";
   IN2_i <= "01010110010001001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100010010";
   IN2_i <= "00010000001010011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101110101";
   IN2_i <= "00011110011101000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111010000";
   IN2_i <= "00100010110001010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011111100";
   IN2_i <= "00000101101000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001110111";
   IN2_i <= "01100000010000000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111101";
   IN2_i <= "01011100110100101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000100110";
   IN2_i <= "01101100110010101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011111010";
   IN2_i <= "00110000000101010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000100000";
   IN2_i <= "00001100010101001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110110111";
   IN2_i <= "00100011000010010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101001111";
   IN2_i <= "01110000101000100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010100100";
   IN2_i <= "00010100111010110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011010110";
   IN2_i <= "00100100011100110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110001001";
   IN2_i <= "00010010100111101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111000100";
   IN2_i <= "00100111001100101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001000100";
   IN2_i <= "01111010011010101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010001101";
   IN2_i <= "00011011010101110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110111101";
   IN2_i <= "00101101110100100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000010111";
   IN2_i <= "00001001001000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110001100";
   IN2_i <= "01010111110110100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111001000";
   IN2_i <= "00001101110110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101100001";
   IN2_i <= "01101000001110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111011111";
   IN2_i <= "01000110100110110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010100";
   IN2_i <= "00100100100101111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100000110";
   IN2_i <= "01100001110101111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101101010";
   IN2_i <= "01010011100100101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110111100";
   IN2_i <= "01001111011010000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000010000";
   IN2_i <= "01011010100110010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101001111";
   IN2_i <= "01001000011011011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100110000";
   IN2_i <= "00100100111101001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010000101";
   IN2_i <= "01000010000000011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100011011";
   IN2_i <= "00011111110010101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010011100";
   IN2_i <= "01101000100010001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011111";
   IN2_i <= "01000000100110111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100000001";
   IN2_i <= "01100011001101010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001111100";
   IN2_i <= "01101100001100101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101011110";
   IN2_i <= "00010010101110000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111101000";
   IN2_i <= "01000010101110011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001100000";
   IN2_i <= "01111011001010110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110110100";
   IN2_i <= "00011100110011010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110111100";
   IN2_i <= "01111001101010110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100011101";
   IN2_i <= "00011000111000000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111100111";
   IN2_i <= "00101100110100000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010000000";
   IN2_i <= "00000001111000001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110100010";
   IN2_i <= "01010111111011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010101";
   IN2_i <= "00001110001111110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100011110";
   IN2_i <= "00110101110100111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110111111";
   IN2_i <= "00101111111001000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100111";
   IN2_i <= "01110001000101011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110101000";
   IN2_i <= "01000110101100110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101000001";
   IN2_i <= "00101011000000010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111011010";
   IN2_i <= "01000001101011111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010100011";
   IN2_i <= "01010000111100101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001110101";
   IN2_i <= "00001100101100110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010100000";
   IN2_i <= "01110010011100001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110001";
   IN2_i <= "00011111001111010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001010111";
   IN2_i <= "00100111001101011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110011110";
   IN2_i <= "00111010010001001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010000010";
   IN2_i <= "01111010111100111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000000011";
   IN2_i <= "01110010010011010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110011001";
   IN2_i <= "00101111000111001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000111011";
   IN2_i <= "01000011011101011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111101101";
   IN2_i <= "01011010110011000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011011111";
   IN2_i <= "00000001000111010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000101011";
   IN2_i <= "01000011010001011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010100111";
   IN2_i <= "01101111101100101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110100000";
   IN2_i <= "01101010111010000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001101011";
   IN2_i <= "01000111110100101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011101011";
   IN2_i <= "01110100110111111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100011011";
   IN2_i <= "01100000100111000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110001000";
   IN2_i <= "01001101100010000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110100101";
   IN2_i <= "01010111100100011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100000111";
   IN2_i <= "00001110100110001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011010000";
   IN2_i <= "01011101101011000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111100010";
   IN2_i <= "00001000011001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100010111";
   IN2_i <= "01100111100100110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000000111";
   IN2_i <= "00000010100010000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011000111";
   IN2_i <= "00011110010011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011000111";
   IN2_i <= "00110011111100110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110000110";
   IN2_i <= "01100100000011101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110101010";
   IN2_i <= "00011111100101011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010001010";
   IN2_i <= "01101011010000001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100011111";
   IN2_i <= "00110001101011001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010101";
   IN2_i <= "00011010011100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011111110";
   IN2_i <= "01000110010100110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100101011";
   IN2_i <= "00111011111010100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000000110";
   IN2_i <= "00000001001001101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010010101";
   IN2_i <= "01111001000010101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000000110";
   IN2_i <= "00110001010110111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011001101";
   IN2_i <= "01011001101001101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000111110";
   IN2_i <= "01101010101100111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100000010";
   IN2_i <= "00001100001001100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111010001";
   IN2_i <= "00101011111011001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101000001";
   IN2_i <= "01100010011100000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101101111";
   IN2_i <= "00010001110011000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100000010";
   IN2_i <= "00101110000100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101000011";
   IN2_i <= "01010101111100010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100001111";
   IN2_i <= "00000111100001101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010110011";
   IN2_i <= "00010100111111111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100011010";
   IN2_i <= "00001101001101100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111011001";
   IN2_i <= "00000110101110001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101101001";
   IN2_i <= "01110010011000000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101100";
   IN2_i <= "00100101110111111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011101000";
   IN2_i <= "01100000010000011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010111101";
   IN2_i <= "00000011100001100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111111111";
   IN2_i <= "01110111101111110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000011100";
   IN2_i <= "00110101011100000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001011110";
   IN2_i <= "00000000100101100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110011001";
   IN2_i <= "01000010100110001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010000";
   IN2_i <= "01001001111011111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101000101";
   IN2_i <= "01101010111110101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000000";
   IN2_i <= "01111100100110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011111001";
   IN2_i <= "00000001011111101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101011101";
   IN2_i <= "01110011011101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001111111";
   IN2_i <= "00100101110010011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110010011";
   IN2_i <= "00011101010000100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111101000";
   IN2_i <= "01111001000111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001011011";
   IN2_i <= "00011100010010100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010011011";
   IN2_i <= "01101001101010000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010101000";
   IN2_i <= "00011111110011001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011101101";
   IN2_i <= "00111100101100101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101000101";
   IN2_i <= "01000010100010100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001010000";
   IN2_i <= "01011010101011101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100110001";
   IN2_i <= "01011100100110101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111101010";
   IN2_i <= "01000011111011011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011000011";
   IN2_i <= "01110011010101101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011111011";
   IN2_i <= "00111100110000110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000110110";
   IN2_i <= "01110111111110010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110000100";
   IN2_i <= "00001111000000101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100010111";
   IN2_i <= "00000010110001100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101001100";
   IN2_i <= "01101101111111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101111011";
   IN2_i <= "00001010110101110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011100100";
   IN2_i <= "01101001101001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101011010";
   IN2_i <= "01110001101111001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111101";
   IN2_i <= "01001011000000011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001010100";
   IN2_i <= "00000010100111001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000101101";
   IN2_i <= "00111100010000010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010010110";
   IN2_i <= "00101001000111011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111011010";
   IN2_i <= "00001100010100110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100100001";
   IN2_i <= "00110000001100100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101000100";
   IN2_i <= "00011001111111110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011001110";
   IN2_i <= "01010111001100000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111001100";
   IN2_i <= "01100001111001111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001110111";
   IN2_i <= "01011111100010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000110101";
   IN2_i <= "01000111111101001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101100001";
   IN2_i <= "01011110110011010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011001001";
   IN2_i <= "01100010011010010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101110010";
   IN2_i <= "00000100001101000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100011010";
   IN2_i <= "00001100100010111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011101011";
   IN2_i <= "00101100100010101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000111100";
   IN2_i <= "01100100011001111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010000101";
   IN2_i <= "01011110000100110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000101100";
   IN2_i <= "01001011101000100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101100011";
   IN2_i <= "00100101010001110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111101110";
   IN2_i <= "00010010101111011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000101011";
   IN2_i <= "00101000010100100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100100001";
   IN2_i <= "00111101100101101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010101111";
   IN2_i <= "01001101000001100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101101101";
   IN2_i <= "01111010100110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100100000";
   IN2_i <= "00011101011101110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011001110";
   IN2_i <= "01101001011111101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110010010";
   IN2_i <= "00110100000000110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001011111";
   IN2_i <= "01100101000000110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110000110";
   IN2_i <= "01011101001100011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001010100";
   IN2_i <= "01010111101001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011101011";
   IN2_i <= "00010101000010011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000100101";
   IN2_i <= "01110001001010100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000011111";
   IN2_i <= "01010010000010010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010100000";
   IN2_i <= "01000000001000111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101011011";
   IN2_i <= "00111110100100010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011100010";
   IN2_i <= "01101000010100011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000010101";
   IN2_i <= "00000110001111000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011011111";
   IN2_i <= "01100010101000111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011100010";
   IN2_i <= "01010001110100101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101011000";
   IN2_i <= "00011011001100000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011000010";
   IN2_i <= "01110001010111010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111110001";
   IN2_i <= "01010010110001011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000000100";
   IN2_i <= "01100111100000101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100101110";
   IN2_i <= "01101011000111101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101111011";
   IN2_i <= "00101110101110011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111110100";
   IN2_i <= "00110111010110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111101000";
   IN2_i <= "01111100101000111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010001000";
   IN2_i <= "00111001100111010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110100100";
   IN2_i <= "00000110110110000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001010000";
   IN2_i <= "00110010011001110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101100100";
   IN2_i <= "01001111011000001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110100100";
   IN2_i <= "01101101010100100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000011";
   IN2_i <= "01001111100101111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000101";
   IN2_i <= "00101001011111100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010100100";
   IN2_i <= "00000011110101111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111011010";
   IN2_i <= "01010001011001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110000000";
   IN2_i <= "01011111110101111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110011111";
   IN2_i <= "01100001111011011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000101100";
   IN2_i <= "01100000100001110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000100000";
   IN2_i <= "01001101000100011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100110011";
   IN2_i <= "00101101111101000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011010000";
   IN2_i <= "00001011011100100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010100010";
   IN2_i <= "00101101110111100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010101111";
   IN2_i <= "00110101111010011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010111010";
   IN2_i <= "00111001110100100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101011111";
   IN2_i <= "01111001111000111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000011010";
   IN2_i <= "00001000001011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110100110";
   IN2_i <= "01100000010100100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000001000";
   IN2_i <= "00011110101110111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111101000";
   IN2_i <= "01111110111001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011010101";
   IN2_i <= "00001110110101110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010100010";
   IN2_i <= "00101111100100011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110100101";
   IN2_i <= "01110011111101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101010010";
   IN2_i <= "01101000100000101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001000101";
   IN2_i <= "00011110111101110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010011110";
   IN2_i <= "00001000001110000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110100100";
   IN2_i <= "00011101110100111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001110011";
   IN2_i <= "00110011111100011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000010001";
   IN2_i <= "01101001101100100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011010";
   IN2_i <= "01100001111001100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001010100";
   IN2_i <= "01100111110000001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100010011";
   IN2_i <= "01001010110000011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101101";
   IN2_i <= "01010101111111010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110011011";
   IN2_i <= "00010010111101101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011111110";
   IN2_i <= "00111110001010001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101100101";
   IN2_i <= "01001011110000000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001110100";
   IN2_i <= "01101001111001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001010100";
   IN2_i <= "00011111001010001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011011000";
   IN2_i <= "01110100111010101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101000111";
   IN2_i <= "01001010001100110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100100001";
   IN2_i <= "01001001010000001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011011011";
   IN2_i <= "01111000000010010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111100011";
   IN2_i <= "00101110100000001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010001001";
   IN2_i <= "01100111001001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011011010";
   IN2_i <= "00001011010011011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010110";
   IN2_i <= "00101110001010010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001101000";
   IN2_i <= "01000001101011011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111000001";
   IN2_i <= "00110011001110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101111010";
   IN2_i <= "01101100111010101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010011";
   IN2_i <= "01011101111010001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010101";
   IN2_i <= "00111011011001110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011100101";
   IN2_i <= "01100000100101110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010101100";
   IN2_i <= "01110011101011001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110111010";
   IN2_i <= "00101011111100001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001111111";
   IN2_i <= "00000100100011001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110000011";
   IN2_i <= "00101100110111101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101111110";
   IN2_i <= "00110110000100011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101110101";
   IN2_i <= "00011101111011111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011001001";
   IN2_i <= "00001010011100001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111010";
   IN2_i <= "00001010001100100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011000";
   IN2_i <= "01001110111000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011110010";
   IN2_i <= "00001001001010100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111010";
   IN2_i <= "00101001111001011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001000111";
   IN2_i <= "01010110101000010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000101110";
   IN2_i <= "00101011100000001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111010000";
   IN2_i <= "00000000011011011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001001000";
   IN2_i <= "00111101001000101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000000101";
   IN2_i <= "00111101001111010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010011010";
   IN2_i <= "01110000111010000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011110";
   IN2_i <= "00111111011000001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010000000";
   IN2_i <= "00110010011010101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001101011";
   IN2_i <= "01111100100011000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110001100";
   IN2_i <= "00111101111100000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111001111";
   IN2_i <= "01111111111110000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001000011";
   IN2_i <= "01111011011101111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111111101";
   IN2_i <= "00110010111011101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010000011";
   IN2_i <= "01101010100010110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101011011";
   IN2_i <= "01111100001100101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100111111";
   IN2_i <= "01001100100000001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011000000";
   IN2_i <= "00110110110001111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011011001";
   IN2_i <= "01001101110010110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000000";
   IN2_i <= "00101001010101111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011111000";
   IN2_i <= "00010001100101011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011100000";
   IN2_i <= "00111110001001111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111001110";
   IN2_i <= "01100011010101101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100000001";
   IN2_i <= "01000101100011000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011000000";
   IN2_i <= "00010100001110110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111100100";
   IN2_i <= "00001100100011101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000101011";
   IN2_i <= "00110101101101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001001101";
   IN2_i <= "00111011000111101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111111101";
   IN2_i <= "01010011001001011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101110011";
   IN2_i <= "01110011111001000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001111101";
   IN2_i <= "00101011010001101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001011100";
   IN2_i <= "01110000010000100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100101010";
   IN2_i <= "00010111000111110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110010000";
   IN2_i <= "00010110100111011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010000110";
   IN2_i <= "00100010110010110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000100";
   IN2_i <= "01110111111110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000011101";
   IN2_i <= "00111001000100000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111101100";
   IN2_i <= "01001101110001101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010110010";
   IN2_i <= "01101100011011101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101101011";
   IN2_i <= "00011001111111110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000100010";
   IN2_i <= "01011110100111011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011011011";
   IN2_i <= "00000010100110011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100101111";
   IN2_i <= "01111011001000000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010011";
   IN2_i <= "01000001101000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111000001";
   IN2_i <= "01001110011000101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100101001";
   IN2_i <= "01000110110100101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001011001";
   IN2_i <= "00010011110011111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111011011";
   IN2_i <= "01010011101000010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101011101";
   IN2_i <= "01010111101001001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010100101";
   IN2_i <= "01011000100001001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010100010";
   IN2_i <= "01000101111001001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110011100";
   IN2_i <= "00000101010010110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110110101";
   IN2_i <= "00110001111011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000111000";
   IN2_i <= "01010010010111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100000011";
   IN2_i <= "00001110000001010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000101000";
   IN2_i <= "00111111001000010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001011000";
   IN2_i <= "00001101010010001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011100010";
   IN2_i <= "01100110110000010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110101010";
   IN2_i <= "01110010001101010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111001";
   IN2_i <= "01001101110011100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110110001";
   IN2_i <= "00000111000111010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001001001";
   IN2_i <= "01100011111010110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111111011";
   IN2_i <= "00110111111010011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000000101";
   IN2_i <= "01101000010100011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100110110";
   IN2_i <= "01000010001110000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011010111";
   IN2_i <= "00100101100100111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001110110";
   IN2_i <= "00100101010100111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001011001";
   IN2_i <= "01101110101011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101111";
   IN2_i <= "00000111011011110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101001110";
   IN2_i <= "00011001110001111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001001110";
   IN2_i <= "00001000101000000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001010110";
   IN2_i <= "01001101011110111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100110011";
   IN2_i <= "00110100101100110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101100111";
   IN2_i <= "00000110000001100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111100100";
   IN2_i <= "00111001101010101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001011100";
   IN2_i <= "00110010101010000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100111011";
   IN2_i <= "01101010110100011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101010111";
   IN2_i <= "00101101100011001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110011111";
   IN2_i <= "00101110100001000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100000111";
   IN2_i <= "00001111011001001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111101001";
   IN2_i <= "01000010010010100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000010100";
   IN2_i <= "00100010111000001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010101111";
   IN2_i <= "00111111011010100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110011110";
   IN2_i <= "00001110100111101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101011000";
   IN2_i <= "01101101111001010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011010001";
   IN2_i <= "00011010011111001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110010010";
   IN2_i <= "00011001110111110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100011000";
   IN2_i <= "01101011001001101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000100001";
   IN2_i <= "00001100101101101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101000010";
   IN2_i <= "01001011000110110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010011110";
   IN2_i <= "00100111000100011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101111110";
   IN2_i <= "00111100110111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111101110";
   IN2_i <= "00100100110000110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111001101";
   IN2_i <= "01101100111011000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011101111";
   IN2_i <= "01110000000111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001111001";
   IN2_i <= "00000110000111011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101111001";
   IN2_i <= "00001011100011001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101001100";
   IN2_i <= "00111110110001000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001010000";
   IN2_i <= "01110010110100100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001000011";
   IN2_i <= "00011101110111100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001011100";
   IN2_i <= "01110010100111001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000000101";
   IN2_i <= "00100000010110010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100000010";
   IN2_i <= "00000111000111011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100111001";
   IN2_i <= "00110000010101000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110001011";
   IN2_i <= "00010110110100010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101111101";
   IN2_i <= "01101001111110001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001010101";
   IN2_i <= "01101001000111110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010100110";
   IN2_i <= "01000011100001010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110100010";
   IN2_i <= "01010111000111010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010110011";
   IN2_i <= "00010111011110101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110100001";
   IN2_i <= "00111000111011100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110010100";
   IN2_i <= "01101010000001001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100000111";
   IN2_i <= "01100001000100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110101000";
   IN2_i <= "01111100110011111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101110011";
   IN2_i <= "01110001001000010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000000101";
   IN2_i <= "01011111010010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100000";
   IN2_i <= "01011000000111001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010101";
   IN2_i <= "00010011100100001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000100000";
   IN2_i <= "01100101111011011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100111";
   IN2_i <= "00101010001010100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001111010";
   IN2_i <= "00111011101100000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000000001";
   IN2_i <= "01111111101010101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010110";
   IN2_i <= "00010101000111011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001101111";
   IN2_i <= "01010110011111100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111010010";
   IN2_i <= "00110011011011100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010110000";
   IN2_i <= "01010100110010001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001100101";
   IN2_i <= "00100111011111110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110011111";
   IN2_i <= "01101011010100100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001110010";
   IN2_i <= "01011111001100100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010101100";
   IN2_i <= "01010100111100011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111101";
   IN2_i <= "00100111101110011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001101000";
   IN2_i <= "00000010000010111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100000011";
   IN2_i <= "01111101011110101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110001000";
   IN2_i <= "00101011101000101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101000010";
   IN2_i <= "01111010000100100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110010001";
   IN2_i <= "00101000100101101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101011000";
   IN2_i <= "01010100001011000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100101000";
   IN2_i <= "00110111010000111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010110";
   IN2_i <= "00000101100101001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011010";
   IN2_i <= "01110101101100111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011100100";
   IN2_i <= "01011010010011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111011111";
   IN2_i <= "00001101110000011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010010010";
   IN2_i <= "01100100010101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010001001";
   IN2_i <= "01101100110111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111100000";
   IN2_i <= "00000101001100101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110110110";
   IN2_i <= "01111100101100010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111011";
   IN2_i <= "00100110110111101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100001001";
   IN2_i <= "00010100101011001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011100101";
   IN2_i <= "01100000000110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001101110";
   IN2_i <= "00001001110100111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010000010";
   IN2_i <= "01111010001011000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011010100";
   IN2_i <= "00111010011000111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110000010";
   IN2_i <= "00001001000111011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100100010";
   IN2_i <= "00100000001011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101111001";
   IN2_i <= "00101111111010100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010101011";
   IN2_i <= "00010101101001101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101111010";
   IN2_i <= "01111111110101011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100000101";
   IN2_i <= "00101110110111111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011110100";
   IN2_i <= "01110011111001010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110100111";
   IN2_i <= "01101011001010000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000010001";
   IN2_i <= "01011001101001000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011111100";
   IN2_i <= "00111011110001111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000000010";
   IN2_i <= "01110110100100011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010110111";
   IN2_i <= "01001010100111011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010011110";
   IN2_i <= "01000000110110001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111011100";
   IN2_i <= "01111100001001111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010111110";
   IN2_i <= "01101000111000010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011111111";
   IN2_i <= "01100011011110110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100110110";
   IN2_i <= "01111111011110111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101111100";
   IN2_i <= "01001010001010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010111101";
   IN2_i <= "01011101000010110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100011111";
   IN2_i <= "00000010101010010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111010100";
   IN2_i <= "01010100101100100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011100100";
   IN2_i <= "00000001010001101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000001100";
   IN2_i <= "00111000110010101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000000101";
   IN2_i <= "00100000110010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111011010";
   IN2_i <= "00110111001001100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011000001";
   IN2_i <= "00001101111001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011110111";
   IN2_i <= "01001111111011111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001010010";
   IN2_i <= "00011000000111111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110001001";
   IN2_i <= "00001010011111110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010110100";
   IN2_i <= "00100100110001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010010100";
   IN2_i <= "00000110010101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100100";
   IN2_i <= "00100000101111000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001010101";
   IN2_i <= "00001111101010101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110010000";
   IN2_i <= "01100110111010001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001100110";
   IN2_i <= "00101011001110110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101111111";
   IN2_i <= "01011001001011110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001010001";
   IN2_i <= "00110111111100001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011101110";
   IN2_i <= "00000011011010001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101000000";
   IN2_i <= "00011100001001001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001100110";
   IN2_i <= "01011001111010110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100111111";
   IN2_i <= "01110000110111101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111010";
   IN2_i <= "00110010111010100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000001010";
   IN2_i <= "01100111101000100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011010100";
   IN2_i <= "01001010010011111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111100";
   IN2_i <= "00100001110100100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100100";
   IN2_i <= "01001001111000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011000110";
   IN2_i <= "00110010110010001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000010100";
   IN2_i <= "01001100000001011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001110101";
   IN2_i <= "01110011111110101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110101110";
   IN2_i <= "01001011111000100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000001";
   IN2_i <= "01010010010111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011011100";
   IN2_i <= "01001110110110000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011000010";
   IN2_i <= "00111010001101110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100110100";
   IN2_i <= "00001000001010010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111001";
   IN2_i <= "00000001011000010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000010110";
   IN2_i <= "00001001110100001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111100100";
   IN2_i <= "01111110000000111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100100100";
   IN2_i <= "01110010110001011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011010010";
   IN2_i <= "00110011101111010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011101101";
   IN2_i <= "00101011010000111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010000001";
   IN2_i <= "00010010001110011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110001001";
   IN2_i <= "01101010100010100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110000011";
   IN2_i <= "00000011000011000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101000100";
   IN2_i <= "00011101001010011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101111010";
   IN2_i <= "01110010011101111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001111010";
   IN2_i <= "01011100100111110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101001011";
   IN2_i <= "01001010110111011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111011010";
   IN2_i <= "01111001111010100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111111100";
   IN2_i <= "01100111101011111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101111111";
   IN2_i <= "01100010100001001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111010100";
   IN2_i <= "01000111111010011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010000100";
   IN2_i <= "00111000000101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101000001";
   IN2_i <= "01110110000101011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011011111";
   IN2_i <= "01000111100010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110110111";
   IN2_i <= "01011001101000100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100010000";
   IN2_i <= "01010000100011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000010";
   IN2_i <= "00000010110000111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110100100";
   IN2_i <= "01101111010011011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101010010";
   IN2_i <= "00011011111110011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001000011";
   IN2_i <= "01001011101101010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100001110";
   IN2_i <= "00100101100101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000001011";
   IN2_i <= "01111100001111001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111101110";
   IN2_i <= "00101000100011011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110100011";
   IN2_i <= "01000101110110001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100001111";
   IN2_i <= "00010000010001000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011100111";
   IN2_i <= "01011011001001001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000110110";
   IN2_i <= "01011111010011000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110010100";
   IN2_i <= "00010110101111101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011001100";
   IN2_i <= "00100101101111001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000000010";
   IN2_i <= "01100111110010010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111000101";
   IN2_i <= "00100100111111001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100101";
   IN2_i <= "01101000110011010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001101011";
   IN2_i <= "01101001010001001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001000101";
   IN2_i <= "00101001100001100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000111110";
   IN2_i <= "01101110011000000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100010101";
   IN2_i <= "01010111010000000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100111010";
   IN2_i <= "01100111001011100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101101110";
   IN2_i <= "01010101011110100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011100111";
   IN2_i <= "01010101111110011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100100110";
   IN2_i <= "01110000000100110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001100011";
   IN2_i <= "00011100111000010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111011000";
   IN2_i <= "00000010100100111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110110110";
   IN2_i <= "00010010001101001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001010111";
   IN2_i <= "01010111010101110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010100001";
   IN2_i <= "01101100001001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101001";
   IN2_i <= "00100110111101110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000000000";
   IN2_i <= "00100010001111001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000110101";
   IN2_i <= "01100010111001011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100001001";
   IN2_i <= "00011111111011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110000110";
   IN2_i <= "01000110101100100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011011111";
   IN2_i <= "00001000000110101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110010000";
   IN2_i <= "00010101010000110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110101011";
   IN2_i <= "01011011111010110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010101111";
   IN2_i <= "01011001101001100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111000111";
   IN2_i <= "01001100011010011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100001100";
   IN2_i <= "00101101010000100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011001000";
   IN2_i <= "00110001011101010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010000100";
   IN2_i <= "01001010100010100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010011111";
   IN2_i <= "00011000010110110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000111000";
   IN2_i <= "01100110001011010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101110";
   IN2_i <= "00011101000111011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010011";
   IN2_i <= "00101110011110000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100000010";
   IN2_i <= "01111000100001110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111011011";
   IN2_i <= "01011110111011011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110001001";
   IN2_i <= "01011001000101000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100010010";
   IN2_i <= "01100110010111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000100010";
   IN2_i <= "01101110110010101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010101110";
   IN2_i <= "00000000100010110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000110111";
   IN2_i <= "00111100000110101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001100100";
   IN2_i <= "01000111010111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111011";
   IN2_i <= "00101011001100101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100100101";
   IN2_i <= "01110011011110110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100110101";
   IN2_i <= "01101111000000111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001111110";
   IN2_i <= "01100101101111110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011101110";
   IN2_i <= "00001110100010110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100000";
   IN2_i <= "00110000001011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111100001";
   IN2_i <= "00110001000101100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000101010";
   IN2_i <= "01001011110000100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000000111";
   IN2_i <= "00101000101111110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010100111";
   IN2_i <= "00111110001110010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001110011";
   IN2_i <= "00000001111010011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111101001";
   IN2_i <= "00001111000100001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110000000";
   IN2_i <= "00101011101001100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011110101";
   IN2_i <= "01000011011000101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110000011";
   IN2_i <= "00001010001010110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101111001";
   IN2_i <= "01101000011001000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010111111";
   IN2_i <= "01101011110101010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100110010";
   IN2_i <= "00001000010101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101011100";
   IN2_i <= "00010001001001011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001110010";
   IN2_i <= "00111100001101000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011001000";
   IN2_i <= "01111111100001100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000110011";
   IN2_i <= "00000100011110111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011111110";
   IN2_i <= "00100000000101101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110100011";
   IN2_i <= "01001110010111111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110010101";
   IN2_i <= "00011101000010011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111100110";
   IN2_i <= "01111000010011001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000111001";
   IN2_i <= "00010000100001111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101101101";
   IN2_i <= "01101001010000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001011010";
   IN2_i <= "01110010100011101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110011010";
   IN2_i <= "01101010110010101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011100000";
   IN2_i <= "01110110111101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101101010";
   IN2_i <= "00101001011110000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001000000";
   IN2_i <= "01111010111000011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001100010";
   IN2_i <= "00111001011000101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101111000";
   IN2_i <= "01010001111001101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001000";
   IN2_i <= "01010000101111001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101100111";
   IN2_i <= "00001101011111101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011110";
   IN2_i <= "01011001111110111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011011010";
   IN2_i <= "00100101001000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001010110";
   IN2_i <= "01101111101010000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010101001";
   IN2_i <= "00101010101100011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100001010";
   IN2_i <= "01110000101111101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011000100";
   IN2_i <= "01000001101011011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000001";
   IN2_i <= "01010011001100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110100110";
   IN2_i <= "01110111010001011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011010100";
   IN2_i <= "01010000101100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110000";
   IN2_i <= "01111000011110111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101001111";
   IN2_i <= "01100000101000010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100010000";
   IN2_i <= "00001000110001111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010001010";
   IN2_i <= "00111111010000100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101100100";
   IN2_i <= "00001100111111110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100010100";
   IN2_i <= "00010101010111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110111110";
   IN2_i <= "00011111000110000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010110011";
   IN2_i <= "01110010011111100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110110010";
   IN2_i <= "01001010001110100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111011001";
   IN2_i <= "00100111001000100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101010101";
   IN2_i <= "00111110010100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010101010";
   IN2_i <= "00011001111101100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001011001";
   IN2_i <= "00101000101011000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010111110";
   IN2_i <= "00101011111000001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011111100";
   IN2_i <= "00111110101110100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010011010";
   IN2_i <= "01001000111100110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001100110";
   IN2_i <= "00100011010111000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110101001";
   IN2_i <= "00110100111001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110111010";
   IN2_i <= "00011100110101001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010000011";
   IN2_i <= "01010010110111100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010010001";
   IN2_i <= "00111001001000111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000101000";
   IN2_i <= "01100100000011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011110101";
   IN2_i <= "00011111000010000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000011100";
   IN2_i <= "00000011010100001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110011011";
   IN2_i <= "01010110100000010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010001011";
   IN2_i <= "00000111110100011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010111100";
   IN2_i <= "01101101000100110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010001001";
   IN2_i <= "00010101001101111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000110111";
   IN2_i <= "01100000110101110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111010101";
   IN2_i <= "01101101000001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000001";
   IN2_i <= "00100100001101110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100001011";
   IN2_i <= "00010100001010110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110110010";
   IN2_i <= "00000101110001111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010101011";
   IN2_i <= "00010100101110111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001101000";
   IN2_i <= "01000001010110011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000010";
   IN2_i <= "01101010110001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111010110";
   IN2_i <= "01101100011000001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011100111";
   IN2_i <= "00001111010111001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011101111";
   IN2_i <= "00110100010010100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111100110";
   IN2_i <= "01000001111001010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110111011";
   IN2_i <= "00011001001010100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000011";
   IN2_i <= "01011001011000010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100110";
   IN2_i <= "00111101011110100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100001111";
   IN2_i <= "00101100000011110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000010010";
   IN2_i <= "00001011100011111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100000100";
   IN2_i <= "01111110000010101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000111010";
   IN2_i <= "00000010100001000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000101100";
   IN2_i <= "01000011000011010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000000110";
   IN2_i <= "01111000001101111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001001011";
   IN2_i <= "00110100110011011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111010010";
   IN2_i <= "00110001001111101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100010001";
   IN2_i <= "00000111000110100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101000001";
   IN2_i <= "01101001010011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001110000";
   IN2_i <= "01101111010001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101110001";
   IN2_i <= "01010011110001111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010111011";
   IN2_i <= "00100110011011000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010111";
   IN2_i <= "00010100111000110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010101100";
   IN2_i <= "00010000000101100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110011011";
   IN2_i <= "01011000001011000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101111011";
   IN2_i <= "01110101100011011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010100100";
   IN2_i <= "00010101100000011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000000101";
   IN2_i <= "00101110101100000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111101010";
   IN2_i <= "00001101000111010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111110010";
   IN2_i <= "00000101101001100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001101011";
   IN2_i <= "01011000010011000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000000001";
   IN2_i <= "01011000111111101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011100100";
   IN2_i <= "01001010000000111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100011";
   IN2_i <= "01100010010111110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000000";
   IN2_i <= "01000000111111001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101000000";
   IN2_i <= "00001010100000101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111100100";
   IN2_i <= "01011011100000001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011000";
   IN2_i <= "00011100100011101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010011000";
   IN2_i <= "00110000011111100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111001100";
   IN2_i <= "01010101011011000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100010101";
   IN2_i <= "01000000111111100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110110001";
   IN2_i <= "01100000110101000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011010110";
   IN2_i <= "00010011111110000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100010100";
   IN2_i <= "01010001001010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000110";
   IN2_i <= "01100001010011111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011100100";
   IN2_i <= "00111111001110000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000011110";
   IN2_i <= "01101001000110110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001001011";
   IN2_i <= "01111010001101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101001011";
   IN2_i <= "00110001111011000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110000111";
   IN2_i <= "01001001101100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111110001";
   IN2_i <= "00110010000010000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001110010";
   IN2_i <= "00110000011010111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101101101";
   IN2_i <= "01011010011000101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100100010";
   IN2_i <= "00101001111000100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001100000";
   IN2_i <= "00111011010000100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111000011";
   IN2_i <= "00010000000110000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010101000";
   IN2_i <= "00011111011111011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111110001";
   IN2_i <= "01010101000011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010101111";
   IN2_i <= "00111101010101110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000100001";
   IN2_i <= "00000111111000000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110010000";
   IN2_i <= "00010110000110111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101110011";
   IN2_i <= "00100100010000011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010110001";
   IN2_i <= "01011101101101011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010000110";
   IN2_i <= "01000101101100000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011001011";
   IN2_i <= "01101100000000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101010000";
   IN2_i <= "00111100001000101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111011100";
   IN2_i <= "00011100010010001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100010111";
   IN2_i <= "00111101010001111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001100";
   IN2_i <= "01011100110110010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001101011";
   IN2_i <= "01100101000101011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101001010";
   IN2_i <= "00000111111010111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101000000";
   IN2_i <= "00100100100100011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110100010";
   IN2_i <= "00011111111101100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001001001";
   IN2_i <= "00110010001110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100011111";
   IN2_i <= "00100001010001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000101010";
   IN2_i <= "01001111000100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011100101";
   IN2_i <= "01101011010111010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100000000";
   IN2_i <= "01100111010100101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001010";
   IN2_i <= "00001010000100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000100111";
   IN2_i <= "01100110111110010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100110111";
   IN2_i <= "01101000001001001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101110110";
   IN2_i <= "01000000110010011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010001001";
   IN2_i <= "01001100101100110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001000";
   IN2_i <= "00101000000110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011100000";
   IN2_i <= "01111110011010101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000110101";
   IN2_i <= "01011011110000010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100100001";
   IN2_i <= "01010100001111100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000010110";
   IN2_i <= "01010110100010111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010100101";
   IN2_i <= "00011100100111001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001000010";
   IN2_i <= "00001110111110000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001000000";
   IN2_i <= "01000110010011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100000111";
   IN2_i <= "00000010111100111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001110110";
   IN2_i <= "01100101011111100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100010110";
   IN2_i <= "01101110110001010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101110001";
   IN2_i <= "01100000111000001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100111";
   IN2_i <= "00111011010011010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111010101";
   IN2_i <= "01001000101111001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001100";
   IN2_i <= "00010010011010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101011111";
   IN2_i <= "01110011101000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011100100";
   IN2_i <= "01100010100001111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010010";
   IN2_i <= "01100000001000111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100111111";
   IN2_i <= "00010010111001010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101001110";
   IN2_i <= "01000100100000001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101000101";
   IN2_i <= "01101110100010000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110011000";
   IN2_i <= "01011100001100110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011110111";
   IN2_i <= "01111100011100011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110000010";
   IN2_i <= "00001100011011101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101000";
   IN2_i <= "01011010010001010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011111111";
   IN2_i <= "01011110010100001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000100010";
   IN2_i <= "01010100001111111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000011110";
   IN2_i <= "00101110110111111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000101001";
   IN2_i <= "01010000100111010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011100010";
   IN2_i <= "01110111100100000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111111011";
   IN2_i <= "01100010101011111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001101";
   IN2_i <= "00010100011100100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100110111";
   IN2_i <= "01101000110010111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110110010";
   IN2_i <= "00000101100000101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010101111";
   IN2_i <= "00001101111001111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110110001";
   IN2_i <= "01001111100011010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101110010";
   IN2_i <= "01111000000001111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110111110";
   IN2_i <= "01000000010010110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000100110";
   IN2_i <= "00101001001101000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101100101";
   IN2_i <= "00111011111111111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111111000";
   IN2_i <= "00000011001000110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001101100";
   IN2_i <= "00011111000000111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111000";
   IN2_i <= "00000011100101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001000110";
   IN2_i <= "01100101111000000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100011";
   IN2_i <= "00110101011001000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101010110";
   IN2_i <= "00100111111100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010100111";
   IN2_i <= "01010000001101011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100001010";
   IN2_i <= "01000010101110010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100000000";
   IN2_i <= "00000001001010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111001100";
   IN2_i <= "00001101011111010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111000100";
   IN2_i <= "00111000000000100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011000001";
   IN2_i <= "00011100000001110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100010011";
   IN2_i <= "01100001111010000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000110010";
   IN2_i <= "01111001000001011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011100101";
   IN2_i <= "01011101100100101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101111111";
   IN2_i <= "00011010001001011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011100";
   IN2_i <= "01100101101011011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101110";
   IN2_i <= "00010101100100100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110101010";
   IN2_i <= "00110011011101010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111110101";
   IN2_i <= "00001101110101101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111010101";
   IN2_i <= "01000111000101100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101101111";
   IN2_i <= "01111010111110111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000010001";
   IN2_i <= "00000001101011110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100111010";
   IN2_i <= "00011100100110000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101100001";
   IN2_i <= "00101010010000010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101011001";
   IN2_i <= "01010011110110010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101100011";
   IN2_i <= "01110110110011111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100100111";
   IN2_i <= "00111101100000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100000";
   IN2_i <= "01101000000110110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110010011";
   IN2_i <= "00110111001100000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101011000";
   IN2_i <= "01011110101010111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001100010";
   IN2_i <= "00100101101010001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000100000";
   IN2_i <= "01110101000001101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100110111";
   IN2_i <= "00110011000110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100110000";
   IN2_i <= "00110110100111011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000101110";
   IN2_i <= "00111011101110110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111011";
   IN2_i <= "00111111000001111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100001010";
   IN2_i <= "01110010000110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101101000";
   IN2_i <= "00000101101101011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001100111";
   IN2_i <= "00010000000101101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000010000";
   IN2_i <= "00011001001001100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100110011";
   IN2_i <= "00100100110000100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001111100";
   IN2_i <= "00010100000100001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000111110";
   IN2_i <= "01000000001111010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100010011";
   IN2_i <= "01100000000010100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000101";
   IN2_i <= "00000011110100110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011101110";
   IN2_i <= "01110001101111011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000100010";
   IN2_i <= "00111001101011111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001000100";
   IN2_i <= "00000011001011111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011011";
   IN2_i <= "00100011111001110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010000001";
   IN2_i <= "00010011010011101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010000010";
   IN2_i <= "00101101001101100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101010100";
   IN2_i <= "00011000100101000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000111111";
   IN2_i <= "01001011100101101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000001001";
   IN2_i <= "00110110000100010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001111110";
   IN2_i <= "00010000100100000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001100101";
   IN2_i <= "01110110011000101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000010101";
   IN2_i <= "01011010101011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100100";
   IN2_i <= "01010010000010010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101011000";
   IN2_i <= "01110111010001101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111101011";
   IN2_i <= "00100110010011101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101001011";
   IN2_i <= "01001000011000110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011101100";
   IN2_i <= "00011100110011110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010011001";
   IN2_i <= "00100111000000110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010101011";
   IN2_i <= "01001001100110010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100110010";
   IN2_i <= "01100000101010010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110110001";
   IN2_i <= "01011001001101011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111001110";
   IN2_i <= "00001101011001101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000011100";
   IN2_i <= "00101111001111001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100100111";
   IN2_i <= "01001111011001000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010001101";
   IN2_i <= "00111111101110101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100111";
   IN2_i <= "00111111010011010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001001111";
   IN2_i <= "00001111011101110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110110111";
   IN2_i <= "01100101011100001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011000110";
   IN2_i <= "00111100000110100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111101001";
   IN2_i <= "01101111100101100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001110110";
   IN2_i <= "01011100010000100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011111110";
   IN2_i <= "01101100100001110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010101111";
   IN2_i <= "01000001110100010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111000111";
   IN2_i <= "01011100001001101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110011010";
   IN2_i <= "01100010011001111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111101111";
   IN2_i <= "01001110111101100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101100110";
   IN2_i <= "00101000000000010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001011101";
   IN2_i <= "01001010010100111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110000111";
   IN2_i <= "00010001101011001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100110111";
   IN2_i <= "01111010100011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110110000";
   IN2_i <= "01111110110100111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101101101";
   IN2_i <= "00101010010001011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000011";
   IN2_i <= "01111110011100011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011101100";
   IN2_i <= "01110111100011011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001000101";
   IN2_i <= "00000100001100010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110010000";
   IN2_i <= "01011111011010011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101001011";
   IN2_i <= "00001001010100011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001111011";
   IN2_i <= "01111010111001100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010111010";
   IN2_i <= "00100110010100111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111110111";
   IN2_i <= "01110100111000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001001000";
   IN2_i <= "01001000011010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001101101";
   IN2_i <= "00100100011110100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000111010";
   IN2_i <= "00000100100111111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100110100";
   IN2_i <= "01111010110110110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110010101";
   IN2_i <= "00110010000111101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001010";
   IN2_i <= "01001111111001101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011001110";
   IN2_i <= "01111110101110011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101001010";
   IN2_i <= "00110011110010111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110110";
   IN2_i <= "00100001101000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000111101";
   IN2_i <= "01000000011011101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000110000";
   IN2_i <= "01011000100001100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011101110";
   IN2_i <= "01111111110011000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111111010";
   IN2_i <= "01111110010100111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111010100";
   IN2_i <= "00101011000010011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010001100";
   IN2_i <= "01100101100010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111110010";
   IN2_i <= "00111011110000110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000011001";
   IN2_i <= "01010011001010000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101010101";
   IN2_i <= "00110010110010000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100100110";
   IN2_i <= "01001100001000011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101101110";
   IN2_i <= "00101011111001110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110111000";
   IN2_i <= "00001110001011100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000001000";
   IN2_i <= "01111011110001000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110111";
   IN2_i <= "00001011101011100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001101011";
   IN2_i <= "00101011011101110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001101001";
   IN2_i <= "00011110101011110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001111111";
   IN2_i <= "00011000110101101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101000111";
   IN2_i <= "00000100000001000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001000100";
   IN2_i <= "01011100110000110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010000011";
   IN2_i <= "00111011010010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011001110";
   IN2_i <= "00100110100001101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011110000";
   IN2_i <= "01101110101000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001000001";
   IN2_i <= "00010011001000000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111000100";
   IN2_i <= "00110110110111110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101011110";
   IN2_i <= "00000111011111110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000010101";
   IN2_i <= "00000100001110011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100100101";
   IN2_i <= "00110011001101111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010011";
   IN2_i <= "01000111000100001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110100100";
   IN2_i <= "01011111010100001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001000001";
   IN2_i <= "00111100000100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001101111";
   IN2_i <= "01010100001100001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000110010";
   IN2_i <= "00110011001100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111001001";
   IN2_i <= "01101010111101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100100";
   IN2_i <= "01001010001010100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010010011";
   IN2_i <= "01011001011101001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111001111";
   IN2_i <= "00001101000101100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101110";
   IN2_i <= "01001011111110111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000110011";
   IN2_i <= "01001101011110010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110111000";
   IN2_i <= "00101100001011010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100010011";
   IN2_i <= "01001010111100100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110010110";
   IN2_i <= "00010011010010110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101011010";
   IN2_i <= "00000011011110111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111010111";
   IN2_i <= "01001000001111000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110110011";
   IN2_i <= "00001011111011100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010010110";
   IN2_i <= "00011110001001000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111111110";
   IN2_i <= "01100111010100000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010011101";
   IN2_i <= "00010110100101010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101001101";
   IN2_i <= "00100011001111111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000000100";
   IN2_i <= "00001000000001101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100000001";
   IN2_i <= "01010001101011110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010101101";
   IN2_i <= "01100001001110001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100100000";
   IN2_i <= "00001010111110001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010010001";
   IN2_i <= "01000000011011100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001101001";
   IN2_i <= "00101101100000101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000001101";
   IN2_i <= "01100111101110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011100111";
   IN2_i <= "00011000100000001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110111000";
   IN2_i <= "00010000000011001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011011001";
   IN2_i <= "01111010111001101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110110010";
   IN2_i <= "01001100010011100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000000010";
   IN2_i <= "00101111110101010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100001110";
   IN2_i <= "00010101100000100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001011101";
   IN2_i <= "00100000001111101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001100001";
   IN2_i <= "00110001010001010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011011101";
   IN2_i <= "00101111000111011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111011";
   IN2_i <= "01100010011111101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000101110";
   IN2_i <= "01000010111100011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000010000";
   IN2_i <= "00111010000001001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011111101";
   IN2_i <= "00101010001000111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011011000";
   IN2_i <= "01100100101101011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101100010";
   IN2_i <= "01110111011111010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010011110";
   IN2_i <= "00110000100100101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010001111";
   IN2_i <= "00101111110011001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111001101";
   IN2_i <= "00000110101101000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001101101";
   IN2_i <= "01000110111001000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001110011";
   IN2_i <= "01111111110010000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111011010";
   IN2_i <= "00010101000010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101001101";
   IN2_i <= "01111110100001100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000010100";
   IN2_i <= "00100011101001010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010010110";
   IN2_i <= "01100010000000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110110111";
   IN2_i <= "01001000011000001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011001011";
   IN2_i <= "01011110110101100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110100010";
   IN2_i <= "01011100001001100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001100010";
   IN2_i <= "01101011110110100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000110100";
   IN2_i <= "01101000011000010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000101";
   IN2_i <= "00111001011010111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101000110";
   IN2_i <= "01110101000111110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001101001";
   IN2_i <= "00111100110001010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110011001";
   IN2_i <= "00100111101110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010101000";
   IN2_i <= "01101011000101100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011010111";
   IN2_i <= "00111100110011001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000010111";
   IN2_i <= "01001001010101011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111101110";
   IN2_i <= "01000110010100101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100111100";
   IN2_i <= "01101110111110111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110110";
   IN2_i <= "00011011111010010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110011010";
   IN2_i <= "01100110100101110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111110000";
   IN2_i <= "01111100000111111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011000101";
   IN2_i <= "01111101000111001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001100111";
   IN2_i <= "00111100111110011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111000";
   IN2_i <= "00110101010001001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101101011";
   IN2_i <= "00000000100110011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100010010";
   IN2_i <= "00010101101110111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111111111";
   IN2_i <= "00101110111000000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110100000";
   IN2_i <= "00011010100110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100000100";
   IN2_i <= "00010011111101100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011100111";
   IN2_i <= "00010001110101001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100001101";
   IN2_i <= "00011100100011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110000011";
   IN2_i <= "01111001101111011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110110001";
   IN2_i <= "01011000011011001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111010011";
   IN2_i <= "01011011001101111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010011001";
   IN2_i <= "01010010001111000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011110010";
   IN2_i <= "00001100000101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001011111";
   IN2_i <= "00110111001000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001101";
   IN2_i <= "00101101001001110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000110110";
   IN2_i <= "00001011110001101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000100011";
   IN2_i <= "01001101010111111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010100100";
   IN2_i <= "01101110010000100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100010011";
   IN2_i <= "00001011000101101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110100001";
   IN2_i <= "01101001101110100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101101010";
   IN2_i <= "00110000011110111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011100010";
   IN2_i <= "01111011010101011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011111";
   IN2_i <= "00011001010011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010000010";
   IN2_i <= "00000010000000000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100000001";
   IN2_i <= "01011010000001111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110111110";
   IN2_i <= "00111101110110111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000001100";
   IN2_i <= "00010001000011100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000100";
   IN2_i <= "00000001110100111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101001010";
   IN2_i <= "01001010011101100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011111010";
   IN2_i <= "01000100011110011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000011000";
   IN2_i <= "01011100010001101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001100100";
   IN2_i <= "00011001011100101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000001101";
   IN2_i <= "01000000011100111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011110";
   IN2_i <= "00100110101011001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100110111";
   IN2_i <= "01000010011110111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001011100";
   IN2_i <= "01001100110000100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001010101";
   IN2_i <= "00011000100111101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010101010";
   IN2_i <= "01110100101000000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010010100";
   IN2_i <= "01011100100101100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111110000";
   IN2_i <= "00110001110101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011101011";
   IN2_i <= "00110010110001110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011101000";
   IN2_i <= "01111110011010001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110011";
   IN2_i <= "01101001011111001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101101111";
   IN2_i <= "01101110010010001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100110";
   IN2_i <= "01001101100100111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101101111";
   IN2_i <= "01001011110000101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011001110";
   IN2_i <= "01100111000111011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101110110";
   IN2_i <= "00001111110011000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001101111";
   IN2_i <= "01001111011001000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000001";
   IN2_i <= "00001011001100101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111111001";
   IN2_i <= "00100100000100001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110101010";
   IN2_i <= "00111011000100111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001110";
   IN2_i <= "01001011101111110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001010011";
   IN2_i <= "00111101001101111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110000";
   IN2_i <= "01011110011000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011101100";
   IN2_i <= "00011111001011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111001110";
   IN2_i <= "00000010000100100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101111101";
   IN2_i <= "00111001001000111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000000101";
   IN2_i <= "01100110100011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100111";
   IN2_i <= "00001011000110001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101101101";
   IN2_i <= "01101001111000101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101001010";
   IN2_i <= "01101101010001001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110100000";
   IN2_i <= "00110000000001110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111110000";
   IN2_i <= "01111111001010001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110000010";
   IN2_i <= "01011110010010010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010101110";
   IN2_i <= "00110010111011101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100101001";
   IN2_i <= "01000100101010010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110000011";
   IN2_i <= "00011110001100100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000000001";
   IN2_i <= "01000111101000001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111110011";
   IN2_i <= "01001010110100010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111110100";
   IN2_i <= "01011010000010111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011001010";
   IN2_i <= "01010011101010011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101101110";
   IN2_i <= "01000011101110110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100001011";
   IN2_i <= "00000101101101001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000110111";
   IN2_i <= "00111001011101001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011010010";
   IN2_i <= "01111011001001011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001010011";
   IN2_i <= "00111001010111111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000111010";
   IN2_i <= "01000001011111100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100100000";
   IN2_i <= "01000011011111001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111111100";
   IN2_i <= "01110111111100100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100000011";
   IN2_i <= "00100100110000001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000011100";
   IN2_i <= "01101001000110000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100101";
   IN2_i <= "00011111001110110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101001011";
   IN2_i <= "01101000101001011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101010001";
   IN2_i <= "00001000111111000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110100110";
   IN2_i <= "00000011101000101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001000011";
   IN2_i <= "01111111010110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101110101";
   IN2_i <= "00011010111010111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011011011";
   IN2_i <= "00010000110101111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010011001";
   IN2_i <= "00010101101101000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100101011";
   IN2_i <= "01000011101010111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100001011";
   IN2_i <= "01100100100110101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110101010";
   IN2_i <= "00011010010111001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111011111";
   IN2_i <= "01010101011101011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001000";
   IN2_i <= "01000001101100111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101001100";
   IN2_i <= "01110011001100001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000100";
   IN2_i <= "00100111111001010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100100110";
   IN2_i <= "00000110000000000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010001";
   IN2_i <= "00011100101011010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101001001";
   IN2_i <= "01011100101101011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011001110";
   IN2_i <= "01000001011111010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011100011";
   IN2_i <= "00110111000000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111010000";
   IN2_i <= "01110100111010010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110111010";
   IN2_i <= "00101000000101110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110000000";
   IN2_i <= "01100110010001101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111111000";
   IN2_i <= "00000001010111111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001110";
   IN2_i <= "00000101000010000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000011110";
   IN2_i <= "01101011000110110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001011001";
   IN2_i <= "01110101101101000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010010100";
   IN2_i <= "00110100111110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011100111";
   IN2_i <= "01100001100010100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001111001";
   IN2_i <= "00001100000010101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001101010";
   IN2_i <= "01001000001110000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101110110";
   IN2_i <= "01101000101111100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011101010";
   IN2_i <= "00101101010010011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111000010";
   IN2_i <= "00100011010001010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110111010";
   IN2_i <= "01011110100000000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010101000";
   IN2_i <= "01100100001000000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011000010";
   IN2_i <= "01111001110100111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111101111";
   IN2_i <= "01011100110011000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100000";
   IN2_i <= "00100111100111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110101111";
   IN2_i <= "01110100000111011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101111111";
   IN2_i <= "01011101011001101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110010111";
   IN2_i <= "00100000000011100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110111";
   IN2_i <= "01000111101110101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011101100";
   IN2_i <= "00010111111100111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110110100";
   IN2_i <= "00001000010111111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111001101";
   IN2_i <= "00010100011100010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111110001";
   IN2_i <= "01010110110100101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100010001";
   IN2_i <= "01110010000000101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100010";
   IN2_i <= "01001010010111111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010001001";
   IN2_i <= "01100110001111100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001110110";
   IN2_i <= "00110001101000011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111110011";
   IN2_i <= "01110000101001000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101000010";
   IN2_i <= "01011111001011100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001101010";
   IN2_i <= "00010001010010001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101100100";
   IN2_i <= "00001111100110111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110000101";
   IN2_i <= "01110101011100011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111000001";
   IN2_i <= "01001110111100011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000100111";
   IN2_i <= "00110100111100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111001010";
   IN2_i <= "01000100010111111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010101001";
   IN2_i <= "01110001111101011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010110010";
   IN2_i <= "00001111011101101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001111101";
   IN2_i <= "00110000011110100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100101100";
   IN2_i <= "00010110101100010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000110010";
   IN2_i <= "01111110110110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111001000";
   IN2_i <= "01001001110010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001110100";
   IN2_i <= "00010000101101011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011010000";
   IN2_i <= "00011110010001111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000111000";
   IN2_i <= "00011110110010001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100110111";
   IN2_i <= "01101111001010010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011101";
   IN2_i <= "01010110011111101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110011110";
   IN2_i <= "00110110101110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101101100";
   IN2_i <= "01110000101111100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010111101";
   IN2_i <= "01100000000101100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111110010";
   IN2_i <= "00001110101000000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111100111";
   IN2_i <= "01111011011111111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101110000";
   IN2_i <= "00111001010000001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100101000";
   IN2_i <= "01111001101101000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111101101";
   IN2_i <= "00111100001111101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101011101";
   IN2_i <= "00000010111101000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011010110";
   IN2_i <= "01100100010100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010001100";
   IN2_i <= "00010010111011101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111101";
   IN2_i <= "00010001000000111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001000101";
   IN2_i <= "01000101101100000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011001100";
   IN2_i <= "00011011101001000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110010011";
   IN2_i <= "00011000110001000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101011100";
   IN2_i <= "01101100010011100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000001";
   IN2_i <= "01010100011110111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001100110";
   IN2_i <= "01011100110100111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111101001";
   IN2_i <= "00001000000000010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010011110";
   IN2_i <= "01100101101000110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011010100";
   IN2_i <= "01100000000001000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100010000";
   IN2_i <= "01101001010011001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101010111";
   IN2_i <= "01001011000000011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110110001";
   IN2_i <= "00000000000010101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110110111";
   IN2_i <= "01010101010111010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110100110";
   IN2_i <= "01010011111110000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010100101";
   IN2_i <= "01010110111110111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000111011";
   IN2_i <= "01010101110100000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100011110";
   IN2_i <= "00011010110100110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010100111";
   IN2_i <= "01111100010100010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000110010";
   IN2_i <= "01010000101010001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100100000";
   IN2_i <= "00000010000100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101101100";
   IN2_i <= "00101111100010001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011100011";
   IN2_i <= "01010100010101110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111100111";
   IN2_i <= "00100001100110100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001010011";
   IN2_i <= "00100101111100010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100101100";
   IN2_i <= "00101110000011101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000011111";
   IN2_i <= "01001100001100101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111111001";
   IN2_i <= "00010111111101011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000011110";
   IN2_i <= "01111100010111100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110111001";
   IN2_i <= "00110110010010111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111011010";
   IN2_i <= "01010001111100011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100101000";
   IN2_i <= "01100100010000000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100100110";
   IN2_i <= "00010000001001110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000111101";
   IN2_i <= "00110010010000101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111100001";
   IN2_i <= "01010100001111100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101011111";
   IN2_i <= "00101110001111101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000110";
   IN2_i <= "01010111000110111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000101100";
   IN2_i <= "00111000000111101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100000101";
   IN2_i <= "01101100100110101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000110111";
   IN2_i <= "00001101101100010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100011101";
   IN2_i <= "00010011110111001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010001000";
   IN2_i <= "01011110111111101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101001101";
   IN2_i <= "01011101000100101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111001111";
   IN2_i <= "01000010100001011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011101000";
   IN2_i <= "00110110001110001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101001101";
   IN2_i <= "00100001101100011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011110011";
   IN2_i <= "01010000011001011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100111001";
   IN2_i <= "01000110001011000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010110000";
   IN2_i <= "01101011001011011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010001010";
   IN2_i <= "01110011001100001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000111100";
   IN2_i <= "00010110000000011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010010001";
   IN2_i <= "00111111010111001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101011010";
   IN2_i <= "01010001110001100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011001111";
   IN2_i <= "00101001100110011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010100101";
   IN2_i <= "01101010111111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101101011";
   IN2_i <= "00100010101010101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111011011";
   IN2_i <= "00101101110000100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001110";
   IN2_i <= "00010000011000100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011010101";
   IN2_i <= "01110011011010000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110010010";
   IN2_i <= "00100000100111011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010011101";
   IN2_i <= "01000111011011001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000011111";
   IN2_i <= "01001101000111001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010100011";
   IN2_i <= "01011101111110100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111100111";
   IN2_i <= "01101111110110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111000100";
   IN2_i <= "01010100010111001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100011011";
   IN2_i <= "00010011100000011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011001100";
   IN2_i <= "01000011100110100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001110000";
   IN2_i <= "01010100001101011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001001110";
   IN2_i <= "00100111111101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001100";
   IN2_i <= "00010000100010110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101001010";
   IN2_i <= "00010010001101100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100000010";
   IN2_i <= "01010110000000010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001110111";
   IN2_i <= "01110110010000100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110000001";
   IN2_i <= "01100100001111111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110001001";
   IN2_i <= "01011101010011100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000100010";
   IN2_i <= "01010010000001010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111100000";
   IN2_i <= "01110100100110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111111000";
   IN2_i <= "00001100110000011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011111101";
   IN2_i <= "01111010111000001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101101100";
   IN2_i <= "01001101001101110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111000101";
   IN2_i <= "01101110101100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110010110";
   IN2_i <= "01110101011100100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010101001";
   IN2_i <= "01110011101110011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000010101";
   IN2_i <= "01110010101010010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100000000";
   IN2_i <= "01111001110101011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111011011";
   IN2_i <= "00111001100010110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111101100";
   IN2_i <= "01101101111100100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000110110";
   IN2_i <= "00110001111110111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011111011";
   IN2_i <= "00110101001111010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000100110";
   IN2_i <= "00100101110010011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001100100";
   IN2_i <= "00001110001100110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011010100";
   IN2_i <= "01111010100110000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001011011";
   IN2_i <= "01100110010100111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101111011";
   IN2_i <= "01000011011010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011101010";
   IN2_i <= "01100011011011000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010101101";
   IN2_i <= "01000101101100101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010010000";
   IN2_i <= "01100111010010000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010010001";
   IN2_i <= "00111110101110100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010100110";
   IN2_i <= "01110010101110000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101010010";
   IN2_i <= "00011011011110000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010001001";
   IN2_i <= "01011001101100101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101100010";
   IN2_i <= "00001011110001001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011011010";
   IN2_i <= "00011001000001110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111000";
   IN2_i <= "01101111011111010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000001000";
   IN2_i <= "01011010011001011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001001000";
   IN2_i <= "01001101001011111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010010";
   IN2_i <= "00000000111101001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111000110";
   IN2_i <= "01001001101100100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100000101";
   IN2_i <= "00010110100011011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110011100";
   IN2_i <= "00111001001000100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010000001";
   IN2_i <= "00110100010110100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110001000";
   IN2_i <= "00001000011010010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111010";
   IN2_i <= "01111100110010010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011010111";
   IN2_i <= "01111101010010100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101000110";
   IN2_i <= "00100000001011100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001001011";
   IN2_i <= "00101111110001011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001110011";
   IN2_i <= "01011010110100100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110110010";
   IN2_i <= "00110010100111001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001111001";
   IN2_i <= "01111110000001010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101101111";
   IN2_i <= "01101111110010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101111010";
   IN2_i <= "00100110010100000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011111101";
   IN2_i <= "01110011000010010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000010000";
   IN2_i <= "00101010100010010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110000001";
   IN2_i <= "01000000101011100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010010111";
   IN2_i <= "01110010100100010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000000000";
   IN2_i <= "01100110001001000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011011000";
   IN2_i <= "01100111100001100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000110000";
   IN2_i <= "01110110101000111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011001001";
   IN2_i <= "00101000000000001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100100010";
   IN2_i <= "01010111011111101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000001111";
   IN2_i <= "01010101001101101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011001100";
   IN2_i <= "00111011101101110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010001111";
   IN2_i <= "00011001100100010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110000011";
   IN2_i <= "00101110001011101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110001101";
   IN2_i <= "01010000010100101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100000000";
   IN2_i <= "01000110001111011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101101011";
   IN2_i <= "01110001000111000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110011001";
   IN2_i <= "00101011011111110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100000";
   IN2_i <= "01110101110011101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000111111";
   IN2_i <= "00111111000011110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110111";
   IN2_i <= "01110111000010011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111110101";
   IN2_i <= "00000000011001000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001010110";
   IN2_i <= "01111110100101100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011000011";
   IN2_i <= "00000111101011010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100011001";
   IN2_i <= "01111010100011000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010111001";
   IN2_i <= "01111111111100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110100100";
   IN2_i <= "01000010011000111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110101101";
   IN2_i <= "01000001000001010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001011";
   IN2_i <= "00000101101011011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000111011";
   IN2_i <= "01111111101000100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100010000";
   IN2_i <= "01001101011100110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101100101";
   IN2_i <= "00110110101101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101111101";
   IN2_i <= "00111010011011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101100011";
   IN2_i <= "00101100001001001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111111010";
   IN2_i <= "00000001011011000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010110100";
   IN2_i <= "00010101110111001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000100100";
   IN2_i <= "01010100011001111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010010110";
   IN2_i <= "01001111111000001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000101010";
   IN2_i <= "00001100110110111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111011000";
   IN2_i <= "01000100010110111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111101";
   IN2_i <= "00110011000010110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001111011";
   IN2_i <= "00101111001100100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111010111";
   IN2_i <= "00101001000100010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000000011";
   IN2_i <= "00011001010101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100001001";
   IN2_i <= "01001110101001100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101101011";
   IN2_i <= "01011101010001000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001100011";
   IN2_i <= "01101100101010011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000110010";
   IN2_i <= "00111100001100100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111100";
   IN2_i <= "00001000010101101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101111010";
   IN2_i <= "00101001011000001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011000010";
   IN2_i <= "00110110000101001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110101010";
   IN2_i <= "00100010101110011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000010001";
   IN2_i <= "00111100110010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011011101";
   IN2_i <= "01000101011111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001010100";
   IN2_i <= "01011011001101001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101010111";
   IN2_i <= "00001101011101110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010010101";
   IN2_i <= "00110101000011001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010011000";
   IN2_i <= "01001000001000010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000100100";
   IN2_i <= "01011011000110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111101";
   IN2_i <= "00011110011100010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111010111";
   IN2_i <= "01101010110100001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100001110";
   IN2_i <= "00010001111100100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000001111";
   IN2_i <= "01100000111101000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001001100";
   IN2_i <= "00100110001010000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110100001";
   IN2_i <= "00000000110100110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010011111";
   IN2_i <= "01000010110010110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000101011";
   IN2_i <= "00011011010001000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011111";
   IN2_i <= "01011011001011101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110010000";
   IN2_i <= "00011110110100000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000000000";
   IN2_i <= "01001010001001001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100010011";
   IN2_i <= "01010111010000111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010011101";
   IN2_i <= "01101100010110001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001011000";
   IN2_i <= "00111101011110110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010010111";
   IN2_i <= "01010010010010000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100111010";
   IN2_i <= "01010100110101000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101100110";
   IN2_i <= "01010011010010110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001111";
   IN2_i <= "00001111101100110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000100110";
   IN2_i <= "01010001011001111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011100100";
   IN2_i <= "00110110111110101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110100111";
   IN2_i <= "00100010111110011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001110101";
   IN2_i <= "00001111111111011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010010010";
   IN2_i <= "00101101100011111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100000010";
   IN2_i <= "01001110001101011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111111001";
   IN2_i <= "00110111101010101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000100001";
   IN2_i <= "01000000001010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101010001";
   IN2_i <= "01110010000110001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101010000";
   IN2_i <= "00011101001001000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111111111";
   IN2_i <= "00100110010001101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110000000";
   IN2_i <= "01000001111011000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100001110";
   IN2_i <= "00010001101000011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101111111";
   IN2_i <= "00000100110101001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101111";
   IN2_i <= "01001101011110001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000001001";
   IN2_i <= "00010011100110110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100110101";
   IN2_i <= "00101010010110010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011110001";
   IN2_i <= "00011110000011110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101001011";
   IN2_i <= "01001111111101101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001101000";
   IN2_i <= "00100011111101001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110100100";
   IN2_i <= "00110001111011100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101010100";
   IN2_i <= "00011010100111010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001011010";
   IN2_i <= "00100001000100011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010110101";
   IN2_i <= "00000010110110001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110011100";
   IN2_i <= "01111111010110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000011010";
   IN2_i <= "01111001000010100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110010";
   IN2_i <= "00111110011001011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111000000";
   IN2_i <= "01000010011000101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000011011";
   IN2_i <= "00000111100100010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011101001";
   IN2_i <= "01100110001110110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000000010";
   IN2_i <= "01100001001110100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111110100";
   IN2_i <= "00010101001001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001100101";
   IN2_i <= "01010100101011111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010000011";
   IN2_i <= "00010100010011100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101001001";
   IN2_i <= "01100001110011101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111011111";
   IN2_i <= "00010011111000001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100111110";
   IN2_i <= "01000101011000110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010100011";
   IN2_i <= "00100000011001001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101010011";
   IN2_i <= "00111111101101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100100100";
   IN2_i <= "01110100001001110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100101111";
   IN2_i <= "00010111000010101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000011100";
   IN2_i <= "01010011010111101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011100000";
   IN2_i <= "01011010101011001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011111101";
   IN2_i <= "01110101001111110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111001110";
   IN2_i <= "00101000000010011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110100001";
   IN2_i <= "00000100111101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100100100";
   IN2_i <= "01100111001100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000011";
   IN2_i <= "01111010110010010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100011010";
   IN2_i <= "00100101011110100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000110110";
   IN2_i <= "01101110111011011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011001100";
   IN2_i <= "00001011001100101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001010110";
   IN2_i <= "01000010010111111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010000110";
   IN2_i <= "00110001101000011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001110110";
   IN2_i <= "01100011100101101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111100010";
   IN2_i <= "01111000111000010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101000010";
   IN2_i <= "00111001101000001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101011010";
   IN2_i <= "00011100010001100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000100010";
   IN2_i <= "01000000111101111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010111";
   IN2_i <= "01111110111010100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100010011";
   IN2_i <= "00011001111001101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001101000";
   IN2_i <= "01100111000110111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100000011";
   IN2_i <= "01110110011111111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111010101";
   IN2_i <= "01100100111110101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000111001";
   IN2_i <= "00010011010010011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011111011";
   IN2_i <= "01000100100110100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001110";
   IN2_i <= "01000100110010000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100100101";
   IN2_i <= "00001111110111100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100001";
   IN2_i <= "00110010101001111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001001110";
   IN2_i <= "01111000001011010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101100110";
   IN2_i <= "01110110001101011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111110111";
   IN2_i <= "00101100001111010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010101001";
   IN2_i <= "01010101111001001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011011001";
   IN2_i <= "01000000001000010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110110";
   IN2_i <= "00000111000100101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001101101";
   IN2_i <= "00101010011111111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001000001";
   IN2_i <= "00110010111100011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011101011";
   IN2_i <= "01111000011011100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100011101";
   IN2_i <= "01100010001011101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001111110";
   IN2_i <= "00000011100001001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101111000";
   IN2_i <= "00111011101111000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101000001";
   IN2_i <= "00111011101011010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110101111";
   IN2_i <= "00110111001001101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111111001";
   IN2_i <= "00011011101100011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111000100";
   IN2_i <= "01110101110110001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111110010";
   IN2_i <= "01000100100110011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010101000";
   IN2_i <= "00011101100110011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100010110";
   IN2_i <= "00100010010000101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101101010";
   IN2_i <= "00100110101101010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111000000";
   IN2_i <= "00010100111100100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011110010";
   IN2_i <= "00000100001000000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001010";
   IN2_i <= "00110001100011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101100110";
   IN2_i <= "01001011110011100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100001000";
   IN2_i <= "00110111001111001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011110110";
   IN2_i <= "01011110010010000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111011111";
   IN2_i <= "00011010001110001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101000";
   IN2_i <= "01111100111001101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001100111";
   IN2_i <= "00110000100100001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110100010";
   IN2_i <= "01111000110110001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000011010";
   IN2_i <= "01110011110000101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110101111";
   IN2_i <= "01110001001010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111011";
   IN2_i <= "00000010100001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100000001";
   IN2_i <= "01010100011111101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111011010";
   IN2_i <= "01101010000010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001100011";
   IN2_i <= "00000001010001010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001110110";
   IN2_i <= "01110100110100111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100100110";
   IN2_i <= "00100000000101011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001001";
   IN2_i <= "01010101111111111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110000001";
   IN2_i <= "01011100011110110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101100010";
   IN2_i <= "00101101000101000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001011011";
   IN2_i <= "00001000110100011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111100101";
   IN2_i <= "01100011000100001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001011110";
   IN2_i <= "01110001001101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110101010";
   IN2_i <= "00110011011101001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000110110";
   IN2_i <= "00100010011110100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101101000";
   IN2_i <= "01111010000001101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000011100";
   IN2_i <= "00000011010111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110011100";
   IN2_i <= "00001100111110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001100101";
   IN2_i <= "01100001100100010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010000011";
   IN2_i <= "00110011010011111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101011001";
   IN2_i <= "01010100100101010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001110101";
   IN2_i <= "00111110011011100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110001100";
   IN2_i <= "00001100110101100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111111010";
   IN2_i <= "00001101110110111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111010100";
   IN2_i <= "00011111110111010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001110110";
   IN2_i <= "00111000111111101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011110";
   IN2_i <= "00110011111100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101010101";
   IN2_i <= "00110101111101000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100101011";
   IN2_i <= "01000111110101001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001000101";
   IN2_i <= "01111000010111100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000010000";
   IN2_i <= "01011101100010010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001010111";
   IN2_i <= "00011111111100010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001000101";
   IN2_i <= "01101111111110000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110010000";
   IN2_i <= "01010011101010100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001010111";
   IN2_i <= "00101101011010100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110100011";
   IN2_i <= "01001010010010011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000000010";
   IN2_i <= "00100000111011101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100101110";
   IN2_i <= "01001110000010101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010101";
   IN2_i <= "01111010100101000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010001100";
   IN2_i <= "01001010000001000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000011000";
   IN2_i <= "01100010001010100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100110010";
   IN2_i <= "00111101010100000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000010100";
   IN2_i <= "00001101011101100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001101100";
   IN2_i <= "00011111100001100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100000001";
   IN2_i <= "01001100001010001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110001111";
   IN2_i <= "00010010011100000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001101001";
   IN2_i <= "00100001101011011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101100011";
   IN2_i <= "01001001111101001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011000010";
   IN2_i <= "01111110011011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001110111";
   IN2_i <= "01110011110101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001111010";
   IN2_i <= "01111010000000111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111111011";
   IN2_i <= "01000110111000110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100001010";
   IN2_i <= "00101011111110101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000101011";
   IN2_i <= "00011100111011001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011011000";
   IN2_i <= "00101110101011100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001000011";
   IN2_i <= "01101111001111000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011000111";
   IN2_i <= "01111000100111010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011001011";
   IN2_i <= "01110001111010011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011111101";
   IN2_i <= "00110001001100001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101111100";
   IN2_i <= "00010011111011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101101011";
   IN2_i <= "00001000101100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000110010";
   IN2_i <= "00100011101011111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110111100";
   IN2_i <= "01001001010110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110111110";
   IN2_i <= "00100000111010011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111101010";
   IN2_i <= "00010001101101011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011111100";
   IN2_i <= "01100110110110100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100111011";
   IN2_i <= "00101011000101001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000111100";
   IN2_i <= "01010101110110111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001010001";
   IN2_i <= "01000111100111101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100101110";
   IN2_i <= "01001101001110101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110101100";
   IN2_i <= "01010101000110110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001001101";
   IN2_i <= "00100100111011001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010110011";
   IN2_i <= "01100001101001001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001111110";
   IN2_i <= "00010111100011100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111101001";
   IN2_i <= "00111011101000000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101001100";
   IN2_i <= "01110000111100111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101000111";
   IN2_i <= "00101100000110010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000110110";
   IN2_i <= "01000001011110101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100100000";
   IN2_i <= "00011011110101101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000010100";
   IN2_i <= "01010111011001110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110000";
   IN2_i <= "01010110111111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001110001";
   IN2_i <= "00011010011101011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111000011";
   IN2_i <= "00100110111011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011011";
   IN2_i <= "00011011100010001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100100011";
   IN2_i <= "01101111001011111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101010011";
   IN2_i <= "01101001111001000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010011101";
   IN2_i <= "01001001111101110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001100110";
   IN2_i <= "00010000000001101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010011000";
   IN2_i <= "00111011001100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001100011";
   IN2_i <= "00001011110101111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100110";
   IN2_i <= "01011010011010100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001010110";
   IN2_i <= "01101101001111000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101000101";
   IN2_i <= "01110010010110000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000000110";
   IN2_i <= "00111101101000010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001101011";
   IN2_i <= "01011000100011100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011100001";
   IN2_i <= "00010000001111011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111111100";
   IN2_i <= "00101000110000010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010001110";
   IN2_i <= "00100101111100100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110010111";
   IN2_i <= "01101101111010100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011000110";
   IN2_i <= "01100111010001000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010111111";
   IN2_i <= "01001001101111011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000010011";
   IN2_i <= "00010000100000101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000101101";
   IN2_i <= "00001011000000101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000100110";
   IN2_i <= "01010110011101011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100001011";
   IN2_i <= "00101010010000010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110000110";
   IN2_i <= "00001110111001010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101110010";
   IN2_i <= "00101100110111000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001101010";
   IN2_i <= "00110000001011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100100110";
   IN2_i <= "00100001010111110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011011011";
   IN2_i <= "01001110001000010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010100100";
   IN2_i <= "00011010100111000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100110011";
   IN2_i <= "00001110100000110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011101101";
   IN2_i <= "01001011011000010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111101111";
   IN2_i <= "01010001101011111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101111";
   IN2_i <= "01110011000001011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111000010";
   IN2_i <= "01110110101101010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110101100";
   IN2_i <= "00111011100111011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111100011";
   IN2_i <= "01100100000100100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000000001";
   IN2_i <= "01101110100110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100000001";
   IN2_i <= "00000100111111010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001011001";
   IN2_i <= "01100001001000101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100000";
   IN2_i <= "00001111101010111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011011111";
   IN2_i <= "01010001011000000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100010110";
   IN2_i <= "01100110111111000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101001110";
   IN2_i <= "01001111010101011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000101110";
   IN2_i <= "00111011000101110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011110000";
   IN2_i <= "00111110011010000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011011010";
   IN2_i <= "00011101100111111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101101001";
   IN2_i <= "01011110011101001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110010010";
   IN2_i <= "01100110010101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100110100";
   IN2_i <= "01001100010111001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000000000";
   IN2_i <= "01000101001011100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011100011";
   IN2_i <= "01101101111110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011010111";
   IN2_i <= "01100001000001001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001010011";
   IN2_i <= "01011010010000011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011111101";
   IN2_i <= "00110111010100101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110101101";
   IN2_i <= "00111000111000010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001010001";
   IN2_i <= "00110011000001100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100110111";
   IN2_i <= "00001011001100100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101011011";
   IN2_i <= "01111010010101110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101101011";
   IN2_i <= "00011011100011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011011010";
   IN2_i <= "00101011101001010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111000";
   IN2_i <= "00001000001000000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111010011";
   IN2_i <= "00100111110111010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010010";
   IN2_i <= "00111101010100111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110011111";
   IN2_i <= "00011111001111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010000101";
   IN2_i <= "00111000010000000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001101100";
   IN2_i <= "01011010101100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101000110";
   IN2_i <= "00001111100011100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001000011";
   IN2_i <= "01010101001100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001010101";
   IN2_i <= "00010110011000101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000000100";
   IN2_i <= "00101101010111010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111100101";
   IN2_i <= "01111101010101110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100110010";
   IN2_i <= "01101010010000110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011001100";
   IN2_i <= "01100001111101101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110011101";
   IN2_i <= "00100110110011011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111011110";
   IN2_i <= "01011001101110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100100111";
   IN2_i <= "00001000101101001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110100001";
   IN2_i <= "01101111101111011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001010101";
   IN2_i <= "00101101100100010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000110111";
   IN2_i <= "00111111101100000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000111101";
   IN2_i <= "01000001000100001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010010011";
   IN2_i <= "01000101101010110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100101110";
   IN2_i <= "00110111100000111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101111011";
   IN2_i <= "00010001011000000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111101101";
   IN2_i <= "00000101011000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010101100";
   IN2_i <= "00111000001001101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011101100";
   IN2_i <= "01110000111110001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001011000";
   IN2_i <= "00000110111110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010101";
   IN2_i <= "00010010100000011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111001";
   IN2_i <= "01111110011000110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011000111";
   IN2_i <= "01010001011110101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010110101";
   IN2_i <= "01000110101100100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011100000";
   IN2_i <= "00110011111000011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010001010";
   IN2_i <= "01111111011010100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010101101";
   IN2_i <= "01101011100101111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101101010";
   IN2_i <= "00110000100100001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100010";
   IN2_i <= "01010100000001100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110011011";
   IN2_i <= "01000010010101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001110101";
   IN2_i <= "00110000101010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111001110";
   IN2_i <= "01111011100000110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001101110";
   IN2_i <= "00101011110011101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101111000";
   IN2_i <= "00111110101010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010110000";
   IN2_i <= "00011100001011000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111011001";
   IN2_i <= "00110001011100101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001001100";
   IN2_i <= "01111001100010101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010010";
   IN2_i <= "01110001010010100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010100000";
   IN2_i <= "01011110001000000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001101";
   IN2_i <= "00000001100000011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010011111";
   IN2_i <= "01000101110100010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100101011";
   IN2_i <= "01110010101111010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101010";
   IN2_i <= "01111101110101101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100000";
   IN2_i <= "00101110000111011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000001100";
   IN2_i <= "00100000110101001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111000111";
   IN2_i <= "00111101101110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100011";
   IN2_i <= "01000001001010101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010110100";
   IN2_i <= "01101000101100001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011101101";
   IN2_i <= "01100101101111010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000010111";
   IN2_i <= "01100000011001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110101101";
   IN2_i <= "00100110001110001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100011000";
   IN2_i <= "00011110111000101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000100000";
   IN2_i <= "01101110011011011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001010101";
   IN2_i <= "01000010001000110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111110011";
   IN2_i <= "00101001111001010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110000011";
   IN2_i <= "01111111010010110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101000001";
   IN2_i <= "00110110001011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010010";
   IN2_i <= "00001010111000110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001101001";
   IN2_i <= "01011010101100011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110010001";
   IN2_i <= "00110011110000001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000100011";
   IN2_i <= "00000001110001110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101111100";
   IN2_i <= "00010101001001111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011111001";
   IN2_i <= "01110110100101100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010110101";
   IN2_i <= "00100101100100001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110001111";
   IN2_i <= "01010000011110101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111110111";
   IN2_i <= "00110011110000101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100010000";
   IN2_i <= "00110111010001110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001000111";
   IN2_i <= "01111100001000101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101011100";
   IN2_i <= "01101111010011000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111101100";
   IN2_i <= "01001100001010111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101101110";
   IN2_i <= "00001110101101001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101001001";
   IN2_i <= "01000100111011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110001111";
   IN2_i <= "00111000011100001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110110011";
   IN2_i <= "00010101000110010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011111000";
   IN2_i <= "00011100011110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001110001";
   IN2_i <= "00010101100110011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001001101";
   IN2_i <= "01100011011000100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010010000";
   IN2_i <= "01110110011110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010000011";
   IN2_i <= "01011010011001101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101111101";
   IN2_i <= "01100011011010101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100010";
   IN2_i <= "00100110000010000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101100100";
   IN2_i <= "00001011011101010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010000101";
   IN2_i <= "00001110100111110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101110101";
   IN2_i <= "00111010000100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101110";
   IN2_i <= "01000010011000101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000101000";
   IN2_i <= "00010000100001101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110101100";
   IN2_i <= "01111101111001100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000010101";
   IN2_i <= "01011000111000100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100101010";
   IN2_i <= "00101010110111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011001000";
   IN2_i <= "00011010110000110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010101101";
   IN2_i <= "00011111100111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111100111";
   IN2_i <= "01110100111000100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110101101";
   IN2_i <= "01011000100011111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100110001";
   IN2_i <= "01000100111111010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101100001";
   IN2_i <= "00010011101111100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101010010";
   IN2_i <= "01001001001010101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100111110";
   IN2_i <= "00010001100010100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010111111";
   IN2_i <= "01011111100100101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000111";
   IN2_i <= "00111000100111110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000110";
   IN2_i <= "01110010011000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110001001";
   IN2_i <= "00010011001111111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100110000";
   IN2_i <= "01010000001111100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010100001";
   IN2_i <= "01111110000011010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110100011";
   IN2_i <= "00010001001111110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001111100";
   IN2_i <= "01101101010100111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000000011";
   IN2_i <= "01101111101101111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111100110";
   IN2_i <= "00110000001001010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111100011";
   IN2_i <= "01110111110000110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000110000";
   IN2_i <= "01001011001100100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010110001";
   IN2_i <= "01000110011101111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001001010";
   IN2_i <= "01101010101011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001000001";
   IN2_i <= "01110101110010111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100011";
   IN2_i <= "01111101101101100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110000000";
   IN2_i <= "01110011110100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001101";
   IN2_i <= "00000101101010011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011110001";
   IN2_i <= "01011000101001100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001001010";
   IN2_i <= "01110101011100000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000110100";
   IN2_i <= "01111000111100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110100011";
   IN2_i <= "00000101010110000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100110000";
   IN2_i <= "00111101101000011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101101";
   IN2_i <= "01001010101001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101100100";
   IN2_i <= "00100010000101001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000011001";
   IN2_i <= "00111110000000111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000101110";
   IN2_i <= "01010001011000100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101010000";
   IN2_i <= "00111010001110101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110000001";
   IN2_i <= "01101001000001110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010010000";
   IN2_i <= "01000100110110011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010001";
   IN2_i <= "01011100010101000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011000101";
   IN2_i <= "01110101010000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111101110";
   IN2_i <= "01010100111011001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101110010";
   IN2_i <= "01100000010011100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110100110";
   IN2_i <= "00110110000010101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100000101";
   IN2_i <= "01000100100001111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101001011";
   IN2_i <= "00011011110100101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001001";
   IN2_i <= "00101011111110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110110010";
   IN2_i <= "00010100011010001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010000001";
   IN2_i <= "00000110100111100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011101111";
   IN2_i <= "01100101110010100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010111101";
   IN2_i <= "00010000010011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100110";
   IN2_i <= "00000010011010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010101000";
   IN2_i <= "00110111001010111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000010011";
   IN2_i <= "00011110101111110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010101010";
   IN2_i <= "01010101100111001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100101000";
   IN2_i <= "00100111001101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000010101";
   IN2_i <= "01101011011101000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101101100";
   IN2_i <= "01101100110011101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110001110";
   IN2_i <= "01011000000111110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100111100";
   IN2_i <= "01001110010111111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100010011";
   IN2_i <= "01011010010101010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000001011";
   IN2_i <= "00101010011000100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001101100";
   IN2_i <= "01011001001000101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110100110";
   IN2_i <= "01101010100111101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110000100";
   IN2_i <= "00010101100000100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010010";
   IN2_i <= "01010001111111011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110010010";
   IN2_i <= "00010111111111101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111001";
   IN2_i <= "01010001010111010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111100100";
   IN2_i <= "00000110100110110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101110101";
   IN2_i <= "00011101011011100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101010110";
   IN2_i <= "01101000001010011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010010101";
   IN2_i <= "01000010100011111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000101111";
   IN2_i <= "01100000001111110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101010";
   IN2_i <= "01001100101111011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010110111";
   IN2_i <= "00111110110010001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001001010";
   IN2_i <= "01101001101000100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100000111";
   IN2_i <= "01101100000001000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000001100";
   IN2_i <= "00000100001101000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101101100";
   IN2_i <= "01001010101110100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100001001";
   IN2_i <= "00110010111100101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101101001";
   IN2_i <= "01100000001010001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100001011";
   IN2_i <= "01010010001011100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010001010";
   IN2_i <= "00111100111101001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000011110";
   IN2_i <= "00001100111001110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111101100";
   IN2_i <= "00101101100011001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001111";
   IN2_i <= "01110001100111110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000011";
   IN2_i <= "01100110100001100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111000111";
   IN2_i <= "00011101110100101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111110001";
   IN2_i <= "00000001100100001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010110110";
   IN2_i <= "01111011011100001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000010110";
   IN2_i <= "01110101010000000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001100";
   IN2_i <= "00011111000110110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110110101";
   IN2_i <= "00010010000100000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001010000";
   IN2_i <= "01110110110111011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110110101";
   IN2_i <= "01111000100111010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100010110";
   IN2_i <= "01110011101001010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110001110";
   IN2_i <= "00001101011011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111111100";
   IN2_i <= "01100011000011001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100010101";
   IN2_i <= "01011001011010011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111010100";
   IN2_i <= "01010110100100011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101110100";
   IN2_i <= "01010100010001110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001011111";
   IN2_i <= "00000010111011000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100110000";
   IN2_i <= "01001110111100000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111001111";
   IN2_i <= "00100111011001110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010100100";
   IN2_i <= "01010000101010110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001000000";
   IN2_i <= "00111100011001111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111100010";
   IN2_i <= "01111110111001000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101101110";
   IN2_i <= "01110111100010110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010101110";
   IN2_i <= "00100001100000100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000100";
   IN2_i <= "01101001110011100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100011100";
   IN2_i <= "00101010000010101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100010";
   IN2_i <= "01001100010111001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100000101";
   IN2_i <= "00111010110101111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011110100";
   IN2_i <= "00111010101000000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011011011";
   IN2_i <= "01010000110111011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000000010";
   IN2_i <= "00011011101111010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111111011";
   IN2_i <= "00001011101100111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101111101";
   IN2_i <= "00110110011111001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110000010";
   IN2_i <= "01010110011001010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000001010";
   IN2_i <= "01111011100010000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001110110";
   IN2_i <= "01001010111111011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001110101";
   IN2_i <= "00010011110101011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100100111";
   IN2_i <= "00011111001100101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101001";
   IN2_i <= "01111000011101111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110101111";
   IN2_i <= "00011111111110000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101010";
   IN2_i <= "01101011000001010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111000111";
   IN2_i <= "00111101010110000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110111110";
   IN2_i <= "00011011001110001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010110010";
   IN2_i <= "00110100111010011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001110101";
   IN2_i <= "00000100000010010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111111010";
   IN2_i <= "00110001110011001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000010110";
   IN2_i <= "01110100001101010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000011111";
   IN2_i <= "01010100011010111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101001001";
   IN2_i <= "00001100100100001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110110011";
   IN2_i <= "00001001100010111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111010111";
   IN2_i <= "01001001001100010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101110010";
   IN2_i <= "01001001001010001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010100010";
   IN2_i <= "01001100011111100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101110001";
   IN2_i <= "00001000010111101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110000100";
   IN2_i <= "00110111011111101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010101";
   IN2_i <= "01010001110101011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111110011";
   IN2_i <= "01000000011011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011100011";
   IN2_i <= "01101100010101011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110000010";
   IN2_i <= "01100000111111001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011011010";
   IN2_i <= "01001000010011011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000001000";
   IN2_i <= "00010000001110001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010110000";
   IN2_i <= "00010111010000100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101001011";
   IN2_i <= "00111100100101111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001111100";
   IN2_i <= "00101011000010000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111000111";
   IN2_i <= "01100010001011111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011111111";
   IN2_i <= "00000010110010000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001111111";
   IN2_i <= "01100000011011101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010101000";
   IN2_i <= "01111111100011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001110011";
   IN2_i <= "01001100111011001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111001111";
   IN2_i <= "01001110101001001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010100011";
   IN2_i <= "00011111111100010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100100001";
   IN2_i <= "01010101000110000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011111010";
   IN2_i <= "01111011011101001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011100110";
   IN2_i <= "00000001011000111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110101000";
   IN2_i <= "01101101010001111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101011101";
   IN2_i <= "00001000010001001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001000110";
   IN2_i <= "01000011100011110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100011011";
   IN2_i <= "00001110100000101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001011100";
   IN2_i <= "00000101001100100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101000011";
   IN2_i <= "00011001001011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000101011";
   IN2_i <= "00111010001001110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011011100";
   IN2_i <= "01110110101001010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000100011";
   IN2_i <= "00010110111101101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001010";
   IN2_i <= "01010010000110001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000111";
   IN2_i <= "00100110110000000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111000100";
   IN2_i <= "00110000111000001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101011";
   IN2_i <= "00001110111111010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110000101";
   IN2_i <= "01011001100110000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111000110";
   IN2_i <= "01101111101001101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111100011";
   IN2_i <= "01101000111101000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100010010";
   IN2_i <= "01101011011100011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101001011";
   IN2_i <= "00011110011110101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100010100";
   IN2_i <= "01011011000010101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011111011";
   IN2_i <= "01111111000111001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001000110";
   IN2_i <= "01100010111010110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011010000";
   IN2_i <= "01101000111010011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001010101";
   IN2_i <= "01110001001110111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001100110";
   IN2_i <= "00010001100000000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111001111";
   IN2_i <= "01001110101011100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111001";
   IN2_i <= "00101111011000101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001110111";
   IN2_i <= "01100000110001011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010110011";
   IN2_i <= "00111101010100011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001011111";
   IN2_i <= "01100100100001001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111101110";
   IN2_i <= "00010110001101100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011101";
   IN2_i <= "01100110001011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111010101";
   IN2_i <= "01010100001101001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001100101";
   IN2_i <= "01100000110000011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001001101";
   IN2_i <= "00100111110100101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101100";
   IN2_i <= "01100110101001110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110000100";
   IN2_i <= "00000011001000001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100000";
   IN2_i <= "00111111010101101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100111";
   IN2_i <= "00101100101111111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001101001";
   IN2_i <= "00010100101001111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110001100";
   IN2_i <= "00101001000100110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101100100";
   IN2_i <= "00010011000100010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000101000";
   IN2_i <= "00101000110001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010101100";
   IN2_i <= "00110010101100100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000011100";
   IN2_i <= "01000011011111010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000110010";
   IN2_i <= "00000100100001111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011100010";
   IN2_i <= "00111001111010101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100111111";
   IN2_i <= "01010110011111011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100011";
   IN2_i <= "01010000110011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001111000";
   IN2_i <= "01100101010011111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111111000";
   IN2_i <= "00111110110100111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100100110";
   IN2_i <= "01111111100010000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111001000";
   IN2_i <= "01101101110100010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001000001";
   IN2_i <= "00000011001001010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001001000";
   IN2_i <= "00111010010110011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100000000";
   IN2_i <= "00010001000101101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011101000";
   IN2_i <= "00101110010111001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011000111";
   IN2_i <= "01110100000100011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101100001";
   IN2_i <= "00110111110010101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000000010";
   IN2_i <= "00101101110001110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101101011";
   IN2_i <= "01001010000001010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100111001";
   IN2_i <= "00101011001000100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100010100";
   IN2_i <= "00010011101100101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110000101";
   IN2_i <= "00101101000001000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111001101";
   IN2_i <= "00101011101111000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111010001";
   IN2_i <= "00011000000100011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100100111";
   IN2_i <= "00110011000100000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010000011";
   IN2_i <= "00110001010100110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100100011";
   IN2_i <= "01000000011000011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100101000";
   IN2_i <= "01101010110111010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010000100";
   IN2_i <= "00010011011000100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010110";
   IN2_i <= "00001011001001101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001101101";
   IN2_i <= "00001101001100100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100100001";
   IN2_i <= "00100111101100110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111111101";
   IN2_i <= "00111000110100000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110100101";
   IN2_i <= "00011100010010111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100101101";
   IN2_i <= "01011010100001100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100001001";
   IN2_i <= "01111101100100010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011010100";
   IN2_i <= "00001101001000101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111011100";
   IN2_i <= "01100101010100001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100101110";
   IN2_i <= "00111010100100110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011100";
   IN2_i <= "01100000100001011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110001010";
   IN2_i <= "01001001001111000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101100010";
   IN2_i <= "00011100011000111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101011000";
   IN2_i <= "00100000100100101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010010";
   IN2_i <= "01110110000011001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001101001";
   IN2_i <= "01110001100000000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110101011";
   IN2_i <= "00000011110101010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000000000";
   IN2_i <= "01100101001100110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011001011";
   IN2_i <= "00011000000000110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010111110";
   IN2_i <= "01100011110110100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000000001";
   IN2_i <= "00110010000001001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000100110";
   IN2_i <= "00101110111001110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110010";
   IN2_i <= "00001001011000110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001000011";
   IN2_i <= "01110100100110110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111110111";
   IN2_i <= "01110000000101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101111001";
   IN2_i <= "01110010100001010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001101000";
   IN2_i <= "00011101010010101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111100111";
   IN2_i <= "00100010111001011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110111000";
   IN2_i <= "00111010100101101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111010111";
   IN2_i <= "01011111011100110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100011101";
   IN2_i <= "01110010000111011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101000110";
   IN2_i <= "00110000110100111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011011100";
   IN2_i <= "00011010111110111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001011110";
   IN2_i <= "00011101110100001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010000011";
   IN2_i <= "01111010001010111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011101011";
   IN2_i <= "01001000010001111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001110110";
   IN2_i <= "01011001000000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011101110";
   IN2_i <= "01100100011011101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100101110";
   IN2_i <= "01110001000001100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010100010";
   IN2_i <= "01100110100110000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010000101";
   IN2_i <= "01001000110011100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011000011";
   IN2_i <= "01101011100000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001110";
   IN2_i <= "01000000000010110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010110111";
   IN2_i <= "01100010111011111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010001001";
   IN2_i <= "01111011001010001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110111";
   IN2_i <= "01001011110110100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101011110";
   IN2_i <= "01110110110110000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100110011";
   IN2_i <= "01101010000111010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100010111";
   IN2_i <= "00111111100111001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111101";
   IN2_i <= "00101001111110011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100110001";
   IN2_i <= "01101000101110100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100000100";
   IN2_i <= "01111010001100101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111001101";
   IN2_i <= "01001100110110101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110011110";
   IN2_i <= "00110100111010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001000000";
   IN2_i <= "01100110001001011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110010111";
   IN2_i <= "00001000011101010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101010010";
   IN2_i <= "00111100100110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100100101";
   IN2_i <= "01100000101110110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000111001";
   IN2_i <= "00110111111111010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101101101";
   IN2_i <= "00011101111000000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100010100";
   IN2_i <= "01001000100110101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000110010";
   IN2_i <= "00101111010000010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011101010";
   IN2_i <= "01000011011000100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101001001";
   IN2_i <= "01011010011111001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101000111";
   IN2_i <= "01000011000111001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010001001";
   IN2_i <= "01101010001010011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111110010";
   IN2_i <= "01011110011111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001001010";
   IN2_i <= "00100101111011100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100110011";
   IN2_i <= "00111100011110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001000101";
   IN2_i <= "01101001001010011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000001011";
   IN2_i <= "00101001010010101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010100100";
   IN2_i <= "01000100101010010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000100001";
   IN2_i <= "01100011110111001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001110101";
   IN2_i <= "00000001110000101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111100001";
   IN2_i <= "01001101100110010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011101001";
   IN2_i <= "00111011110110010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000011101";
   IN2_i <= "01110101011000111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111100011";
   IN2_i <= "01111100100011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011000010";
   IN2_i <= "00001100100010000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101111011";
   IN2_i <= "00101101011011100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101110100";
   IN2_i <= "00010001010101110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101001111";
   IN2_i <= "01001101110111100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100010010";
   IN2_i <= "01011101110101111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000010010";
   IN2_i <= "00100001000001110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100011110";
   IN2_i <= "01001111010000111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101001110";
   IN2_i <= "00010110100001011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001010011";
   IN2_i <= "00101011111101110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111001000";
   IN2_i <= "01001000100001000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100001100";
   IN2_i <= "01000000100110010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111111001";
   IN2_i <= "00110100111111110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001010110";
   IN2_i <= "01001111001001111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001111010";
   IN2_i <= "01000010111011101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101101000";
   IN2_i <= "01001001100110111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111110101";
   IN2_i <= "01110000110111011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110001";
   IN2_i <= "00111011111110000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001100";
   IN2_i <= "00110100001101110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110001000";
   IN2_i <= "01011011111001010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111011010";
   IN2_i <= "01001010100111110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101010110";
   IN2_i <= "00110100100111100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101101";
   IN2_i <= "01000110100100001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001011001";
   IN2_i <= "01100011101010101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011111011";
   IN2_i <= "01101011010101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000000001";
   IN2_i <= "00100111100011100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101110111";
   IN2_i <= "01001001000111100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001011001";
   IN2_i <= "01010101010011011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001010110";
   IN2_i <= "00111100010101010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111101000";
   IN2_i <= "01101010001110110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100001000";
   IN2_i <= "00101110101111111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101101011";
   IN2_i <= "01010101111100101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001000000";
   IN2_i <= "01110100100000001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011110001";
   IN2_i <= "01110111110111100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011110010";
   IN2_i <= "01110001110011111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010100011";
   IN2_i <= "01001010001011001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011010101";
   IN2_i <= "00000111000010000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010001100";
   IN2_i <= "01001000011100100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101010001";
   IN2_i <= "01101100110001010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111101101";
   IN2_i <= "00100001010110001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101101";
   IN2_i <= "00001010111101011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000010011";
   IN2_i <= "01101011100000001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101011100";
   IN2_i <= "01111110000000010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110011001";
   IN2_i <= "00001010001100000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101010000";
   IN2_i <= "01110111101110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110110001";
   IN2_i <= "01110110011011100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001111000";
   IN2_i <= "00001100000001001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000000000";
   IN2_i <= "00010010001010111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101000111";
   IN2_i <= "01000110011101000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111010100";
   IN2_i <= "00110001011100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110011001";
   IN2_i <= "00010000000100100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010011011";
   IN2_i <= "00011000111101110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010111110";
   IN2_i <= "00111001001100111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111100111";
   IN2_i <= "01101110000111101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100111011";
   IN2_i <= "01100110110100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000110100";
   IN2_i <= "01001100101011100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111101011";
   IN2_i <= "00001010111011111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100000011";
   IN2_i <= "00111111110011100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010101010";
   IN2_i <= "01010001010010000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111100";
   IN2_i <= "00111001100100100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011101101";
   IN2_i <= "01100000101001000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101100101";
   IN2_i <= "01010001100000011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001000100";
   IN2_i <= "00110100010110101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100011111";
   IN2_i <= "01111111001010100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100110110";
   IN2_i <= "00001011111001001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110111101";
   IN2_i <= "01010010101110001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000110110";
   IN2_i <= "00100110011001100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100011110";
   IN2_i <= "01100011000000001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010010110";
   IN2_i <= "00101101010010101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011011000";
   IN2_i <= "00111000000010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110011000";
   IN2_i <= "00001010111000110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001011100";
   IN2_i <= "01010011100110001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000010010";
   IN2_i <= "01011001010111100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100011111";
   IN2_i <= "00010000111110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011000111";
   IN2_i <= "00101111001100010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000000";
   IN2_i <= "01111001111010001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110001110";
   IN2_i <= "00100101001101110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111101010";
   IN2_i <= "01101010100110111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100100";
   IN2_i <= "00111010101000100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111000011";
   IN2_i <= "01111010111001100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000110111";
   IN2_i <= "01001110000110010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000111101";
   IN2_i <= "01110100101111011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111000";
   IN2_i <= "01101110011001110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000100101";
   IN2_i <= "00000010110010001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011010010";
   IN2_i <= "01000010110010011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100110000";
   IN2_i <= "01100011101010111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111011010";
   IN2_i <= "00100100101001011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110101001";
   IN2_i <= "00011110110101111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001111";
   IN2_i <= "00111010101011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100100000";
   IN2_i <= "01001011100001101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100011100";
   IN2_i <= "01011110011011011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000100010";
   IN2_i <= "00001100010001010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100110001";
   IN2_i <= "00011110011110110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000001100";
   IN2_i <= "01110010001110110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101001101";
   IN2_i <= "00110101110101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101101100";
   IN2_i <= "01110011011111000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111011101";
   IN2_i <= "01011000100010010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010011101";
   IN2_i <= "00101000011010111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010001001";
   IN2_i <= "01000010100111101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010101110";
   IN2_i <= "01010000011100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001000";
   IN2_i <= "00101110000010010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101001101";
   IN2_i <= "01101101011011011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011101101";
   IN2_i <= "01100001111110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001000";
   IN2_i <= "00110000001011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110010010";
   IN2_i <= "01100100000100110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111100";
   IN2_i <= "01010111110000000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101111100";
   IN2_i <= "00001001001001110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100010100";
   IN2_i <= "01010111001001101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110101000";
   IN2_i <= "01111001011010001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111111011";
   IN2_i <= "00111101111110000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100111010";
   IN2_i <= "00011110111111000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011100111";
   IN2_i <= "00011011110011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110111111";
   IN2_i <= "01000111110000110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101101010";
   IN2_i <= "00010101111111010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001111000";
   IN2_i <= "01000101001011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001010011";
   IN2_i <= "00001001101010110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011111";
   IN2_i <= "00101010110101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100111010";
   IN2_i <= "00011011011001101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111100100";
   IN2_i <= "01000100111001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010100000";
   IN2_i <= "00100010000011101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101001100";
   IN2_i <= "00011111001001110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110101100";
   IN2_i <= "01111111111110001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110001101";
   IN2_i <= "01011010010110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110100101";
   IN2_i <= "00010101011011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111101100";
   IN2_i <= "01111011000010011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000100101";
   IN2_i <= "01100001010001111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110010101";
   IN2_i <= "01000100000110011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111000011";
   IN2_i <= "00111011100010101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101110011";
   IN2_i <= "00111000100100011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110000";
   IN2_i <= "00110000000001011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100010010";
   IN2_i <= "01010010001101100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111001110";
   IN2_i <= "01010100001110000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010001001";
   IN2_i <= "00000110100101100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010011101";
   IN2_i <= "00100011100011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001010000";
   IN2_i <= "00001110101000011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011011000";
   IN2_i <= "00100010001000011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000011000";
   IN2_i <= "01100011110110000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101001111";
   IN2_i <= "01100000100001011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001000";
   IN2_i <= "01100011001111001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001110010";
   IN2_i <= "00100001000001110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010010100";
   IN2_i <= "01011000100011000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000101110";
   IN2_i <= "00111100000010111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010011000";
   IN2_i <= "00001100111010011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010100110";
   IN2_i <= "00100000011000100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101100";
   IN2_i <= "00100101001000011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010010";
   IN2_i <= "00000100000101001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101100111";
   IN2_i <= "01011100110101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101001011";
   IN2_i <= "00110101000000010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100000111";
   IN2_i <= "01011001100110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000110001";
   IN2_i <= "01000110010001010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110010101";
   IN2_i <= "01111111010110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000111011";
   IN2_i <= "00111010010100001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010110";
   IN2_i <= "01100111111110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011000100";
   IN2_i <= "01110110011010010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011000110";
   IN2_i <= "01111110111110101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000110000";
   IN2_i <= "01111111111000111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110001010";
   IN2_i <= "01111110001010000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010000";
   IN2_i <= "01010011011100011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100110101";
   IN2_i <= "00000010000111111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111001010";
   IN2_i <= "00110011100110000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100110011";
   IN2_i <= "01001000001001101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011110101";
   IN2_i <= "01101001000001001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001000110";
   IN2_i <= "01011010101010001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100110100";
   IN2_i <= "00111101111000010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010101110";
   IN2_i <= "00110101100001111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110111011";
   IN2_i <= "00110100010000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010010111";
   IN2_i <= "00010110011001110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110011001";
   IN2_i <= "01110000001001011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001001110";
   IN2_i <= "00110110111111010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101010111";
   IN2_i <= "00010101001000001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101001000";
   IN2_i <= "00011101001011100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011000110";
   IN2_i <= "00111111110001101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011101101";
   IN2_i <= "01011111011011000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111101111";
   IN2_i <= "00101110100101111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101111001";
   IN2_i <= "00100110111101100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011011010";
   IN2_i <= "00011111101000111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010011010";
   IN2_i <= "00101001010001011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100110111";
   IN2_i <= "01111111011110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101110110";
   IN2_i <= "00010111110101011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110110011";
   IN2_i <= "00000101111010100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111011110";
   IN2_i <= "01000110100010110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110101";
   IN2_i <= "01111001111100001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000000111";
   IN2_i <= "00000100000100100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001110001";
   IN2_i <= "01111001100001010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110001110";
   IN2_i <= "01100110011000101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010111011";
   IN2_i <= "01101010000000110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010010000";
   IN2_i <= "00001110101001110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100101001";
   IN2_i <= "00000000011110000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110001";
   IN2_i <= "00100011001110001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010011";
   IN2_i <= "01001011001001100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110001010";
   IN2_i <= "01101110100111010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000001111";
   IN2_i <= "00110100010100100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101010101";
   IN2_i <= "01010110101111100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101111111";
   IN2_i <= "01001111001011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100001100";
   IN2_i <= "00000010010011001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001100";
   IN2_i <= "01011011111100011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011011010";
   IN2_i <= "00110101101001010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001011100";
   IN2_i <= "00101011101010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110111100";
   IN2_i <= "01010110100001000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010111100";
   IN2_i <= "01110100101100000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111001101";
   IN2_i <= "00011010011110100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011110001";
   IN2_i <= "00111011101110110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011101000";
   IN2_i <= "00000111010001001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101101001";
   IN2_i <= "00100011010101010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010111000";
   IN2_i <= "00100011000100101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000111101";
   IN2_i <= "01110010101000010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000101111";
   IN2_i <= "00100011101101010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011110";
   IN2_i <= "00111000010000101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111111";
   IN2_i <= "00011000000001000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111010011";
   IN2_i <= "00100010001110110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001011001";
   IN2_i <= "00101101110010011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111011010";
   IN2_i <= "01101010101111100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100111001";
   IN2_i <= "01100010001110011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001100010";
   IN2_i <= "01110100011010101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001100111";
   IN2_i <= "00001001110011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011001110";
   IN2_i <= "00010011000101010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110011011";
   IN2_i <= "00011000010110011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111100001";
   IN2_i <= "01111111010110110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101101011";
   IN2_i <= "00000010100010110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011011000";
   IN2_i <= "01100110000010001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111100000";
   IN2_i <= "00011010010010011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010001010";
   IN2_i <= "01010110011100001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010001001";
   IN2_i <= "01110001010111001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111101001";
   IN2_i <= "01011011001100101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110010001";
   IN2_i <= "00101011110100111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101100101";
   IN2_i <= "00011101110101101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001111101";
   IN2_i <= "00001000110010111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101010111";
   IN2_i <= "01000110101111110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010011010";
   IN2_i <= "01001111001100010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110011011";
   IN2_i <= "00011111000000011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011000101";
   IN2_i <= "00010110011110100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010100001";
   IN2_i <= "00101110100101101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000001011";
   IN2_i <= "01001110100000011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100000";
   IN2_i <= "01100110000000101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101101100";
   IN2_i <= "00101110100011001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111010010";
   IN2_i <= "01101000110011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001000100";
   IN2_i <= "01110111011100011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101110110";
   IN2_i <= "01011000100001000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100001110";
   IN2_i <= "00001100110111101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010011011";
   IN2_i <= "01000010111010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000100010";
   IN2_i <= "00110010011100101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101100010";
   IN2_i <= "01001000001110010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100110000";
   IN2_i <= "01100011100111000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000100000";
   IN2_i <= "01101100110000011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111100110";
   IN2_i <= "00110011000011110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001110001";
   IN2_i <= "01001011000001101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110000011";
   IN2_i <= "01011100101000100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001010100";
   IN2_i <= "01100000110110100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101010001";
   IN2_i <= "00001100111011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001010011";
   IN2_i <= "01011001111110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111110101";
   IN2_i <= "00010001110101011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101111010";
   IN2_i <= "01001110100100000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001111100";
   IN2_i <= "00111101110100011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010001";
   IN2_i <= "01111110110110001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011001101";
   IN2_i <= "01111000101111111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101100";
   IN2_i <= "01110001101111110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010110011";
   IN2_i <= "01110111010011000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110101010";
   IN2_i <= "01101001111011101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110101";
   IN2_i <= "01111100100110010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110011";
   IN2_i <= "01011100100100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110111001";
   IN2_i <= "01101001001111011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110100";
   IN2_i <= "00010111001100100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001110111";
   IN2_i <= "01001100100100110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011101000";
   IN2_i <= "01010010011101011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101001011";
   IN2_i <= "01000011110011011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001101011";
   IN2_i <= "01010011001011111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100100111";
   IN2_i <= "00101101000011010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001110111";
   IN2_i <= "00110001110010111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011100";
   IN2_i <= "01101001110011010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110010110";
   IN2_i <= "01010000011010001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111100010";
   IN2_i <= "00011110101010100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001001001";
   IN2_i <= "01110111111100010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010100110";
   IN2_i <= "00111010100100110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111111010";
   IN2_i <= "01011100001110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110111100";
   IN2_i <= "00110110101010001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101010010";
   IN2_i <= "01111010010000001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011110000";
   IN2_i <= "00101000110101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100001110";
   IN2_i <= "00010001110110111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101110";
   IN2_i <= "01101000110100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001011010";
   IN2_i <= "01101000110111010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000110000";
   IN2_i <= "00111101110010110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001110000";
   IN2_i <= "00110110010101011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011110100";
   IN2_i <= "00011110011110000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111000000";
   IN2_i <= "01000110101111101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100100110";
   IN2_i <= "01110110101000010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111100101";
   IN2_i <= "01111011010111110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000010000";
   IN2_i <= "00001110111110101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110110000";
   IN2_i <= "00001000011101110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010100000";
   IN2_i <= "01111110011100111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011011101";
   IN2_i <= "00010101110110010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100010110";
   IN2_i <= "00101100110010101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011111101";
   IN2_i <= "00000110001010011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010011101";
   IN2_i <= "01101111110111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110011111";
   IN2_i <= "00110111011111011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000010010";
   IN2_i <= "01011100001011001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001101010";
   IN2_i <= "00101011100101010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111111000";
   IN2_i <= "01101111011010100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001110000";
   IN2_i <= "00010100011011101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011010001";
   IN2_i <= "01011010001100101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110111000";
   IN2_i <= "00001111111011111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000101001";
   IN2_i <= "00101101011110110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000111101";
   IN2_i <= "00100101010000111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000011011";
   IN2_i <= "00100001001000010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001111011";
   IN2_i <= "00110101110111101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110000101";
   IN2_i <= "01000000111011000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110110101";
   IN2_i <= "01100100101110000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111000";
   IN2_i <= "01010111111100100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000011001";
   IN2_i <= "00001010010001111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001010101";
   IN2_i <= "01100010110000001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000101";
   IN2_i <= "01000100111010111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100111111";
   IN2_i <= "00110100110100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000011001";
   IN2_i <= "01010110111011110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011001";
   IN2_i <= "00110011011001011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111010100";
   IN2_i <= "00100011000100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100010101";
   IN2_i <= "00111011100100111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010000001";
   IN2_i <= "01101000000001011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000101";
   IN2_i <= "00110011101001100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000001001";
   IN2_i <= "01011110001010100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111100111";
   IN2_i <= "01000101110001001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011000011";
   IN2_i <= "00001100011001001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011010010";
   IN2_i <= "00011011101111011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001110100";
   IN2_i <= "01100110011101011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100001011";
   IN2_i <= "00111001001011010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100101001";
   IN2_i <= "01000111001001111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111101000";
   IN2_i <= "01010001011110111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010000011";
   IN2_i <= "01101001001100101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100100111";
   IN2_i <= "01101000101011000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101011110";
   IN2_i <= "01001001001010010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001000010";
   IN2_i <= "00111110110110100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110101010";
   IN2_i <= "01101100101010101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001110101";
   IN2_i <= "01101010100000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011000001";
   IN2_i <= "00100000111001111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001011111";
   IN2_i <= "00110111010110101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110001001";
   IN2_i <= "00110001110111101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000110011";
   IN2_i <= "00001011111110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010100011";
   IN2_i <= "00010101101111010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100011";
   IN2_i <= "00101001111110110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010000001";
   IN2_i <= "00011000101000101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111111100";
   IN2_i <= "00001000010000100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100101011";
   IN2_i <= "00110100000001110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010010110";
   IN2_i <= "00100100111111000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100100110";
   IN2_i <= "01010101001111111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100000000";
   IN2_i <= "00101100001010111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100000101";
   IN2_i <= "01010001111000111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010100011";
   IN2_i <= "00011111011000101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010001";
   IN2_i <= "01110011110101010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010100110";
   IN2_i <= "01000100110001111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101000000";
   IN2_i <= "00111110000101000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101101011";
   IN2_i <= "00010111000000001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001100011";
   IN2_i <= "00110100111011001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100101110";
   IN2_i <= "00001110110001100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100101001";
   IN2_i <= "00100001010001100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000111001";
   IN2_i <= "01011000100011011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010110";
   IN2_i <= "00001000001011100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001110101";
   IN2_i <= "01011110010101100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000000011";
   IN2_i <= "01110100001101101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001100010";
   IN2_i <= "01110001011110101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111000001";
   IN2_i <= "01100010100111100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111000101";
   IN2_i <= "00110010010010100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101001011";
   IN2_i <= "01101100011110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101010111";
   IN2_i <= "00111011011101010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110001111";
   IN2_i <= "01011100110001101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111111010";
   IN2_i <= "00010101001001110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110011010";
   IN2_i <= "01011011110110100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001100100";
   IN2_i <= "01111000011010110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110111000";
   IN2_i <= "01000101100101100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001100011";
   IN2_i <= "01001001001101101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000111";
   IN2_i <= "01010101110011010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001111000";
   IN2_i <= "01100101000110100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101000111";
   IN2_i <= "00111111110100011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101010";
   IN2_i <= "00000000000011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000110011000";
   IN2_i <= "01000110100011110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100111";
   IN2_i <= "00011101111010111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101010111";
   IN2_i <= "00000100001011100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001001110";
   IN2_i <= "01110110001010001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111100010";
   IN2_i <= "00000111011010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111110";
   IN2_i <= "01001101101001010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010100111";
   IN2_i <= "01101001101011110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001110";
   IN2_i <= "00110100010100101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110001011";
   IN2_i <= "01010110010010101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010011010";
   IN2_i <= "01101100000101100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000111";
   IN2_i <= "01000110100101000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010110010";
   IN2_i <= "01110001001101010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011111011";
   IN2_i <= "00101101000000010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111000000";
   IN2_i <= "00010101101100100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010110";
   IN2_i <= "00000101110100000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011010110";
   IN2_i <= "01001011101100000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011000011";
   IN2_i <= "00100001010001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101001101";
   IN2_i <= "00000000101111100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111010100";
   IN2_i <= "00000111100000000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000110";
   IN2_i <= "00000100101101000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010011110";
   IN2_i <= "01000110001101101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011100101";
   IN2_i <= "01001001100100101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001110110";
   IN2_i <= "00110010010100100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000011000";
   IN2_i <= "00011111000000011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000011111";
   IN2_i <= "01011000101000001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111010101";
   IN2_i <= "00101111000100111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111011";
   IN2_i <= "01011111000011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011100101";
   IN2_i <= "01010110100100100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101010001";
   IN2_i <= "00011110111001000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000011010";
   IN2_i <= "00111010110101100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011000101";
   IN2_i <= "00011000000111000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110011110";
   IN2_i <= "00011000100000001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000000111";
   IN2_i <= "00010010101001011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101001010";
   IN2_i <= "00110000011111101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011011111";
   IN2_i <= "01100101101100111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101101110";
   IN2_i <= "01010111111111000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001111000";
   IN2_i <= "00011111001100101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000111011";
   IN2_i <= "01001001110011010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000011100";
   IN2_i <= "01000001001101011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101101001";
   IN2_i <= "01011001010010100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011001010";
   IN2_i <= "01001011010101000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011101111";
   IN2_i <= "00101000101111011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110000100";
   IN2_i <= "00110000011100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111111001";
   IN2_i <= "01010011100100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100100100";
   IN2_i <= "00111000101010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000001110";
   IN2_i <= "00010011110001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110100001";
   IN2_i <= "00100100110101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100000000";
   IN2_i <= "00100111110000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000010";
   IN2_i <= "00110011111100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001011010";
   IN2_i <= "01000110011000110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101111001";
   IN2_i <= "01001101011011101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011000011";
   IN2_i <= "01000100000111010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010101111";
   IN2_i <= "00001000110111101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001001011";
   IN2_i <= "01100010011100000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000101010";
   IN2_i <= "01111010101010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101001101";
   IN2_i <= "00011101011100111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010010111";
   IN2_i <= "01111100011001101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001100000";
   IN2_i <= "01101011110000010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111101000";
   IN2_i <= "00110100010111101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011011010";
   IN2_i <= "01110010010110111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101010";
   IN2_i <= "00001100110100111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100100010";
   IN2_i <= "01011101000001100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001110101";
   IN2_i <= "00010111101100010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111111010";
   IN2_i <= "00000110011110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011001011";
   IN2_i <= "01000111100111011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011001010";
   IN2_i <= "01010100010101011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001110";
   IN2_i <= "01100010101101011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011110000";
   IN2_i <= "01110111111011110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000010010";
   IN2_i <= "01011100010100101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010110011";
   IN2_i <= "00011100010010001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001001100";
   IN2_i <= "01011001111110111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100111011";
   IN2_i <= "01101001000000101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010001100";
   IN2_i <= "01101111110100010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000111001";
   IN2_i <= "01110101010111011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010101011";
   IN2_i <= "01100100010101000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000110001";
   IN2_i <= "01101001011011111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111100100";
   IN2_i <= "01100011010110000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100111011";
   IN2_i <= "01010011000001011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111100110";
   IN2_i <= "01011101010011111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010001011";
   IN2_i <= "00101001001000000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010110110";
   IN2_i <= "01011000101110101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001001110";
   IN2_i <= "00011000110011110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011011";
   IN2_i <= "01010100111001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000011010";
   IN2_i <= "00100111010010111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100011100";
   IN2_i <= "00110111010010011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010110011";
   IN2_i <= "00001101010010000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001100011";
   IN2_i <= "00001010000001110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010000100";
   IN2_i <= "01110101000101000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001000";
   IN2_i <= "00101101010011110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111001010";
   IN2_i <= "01111001011000000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101110010";
   IN2_i <= "01111011010000101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100100";
   IN2_i <= "01101000110110001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011110001";
   IN2_i <= "00010111010011000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101110110";
   IN2_i <= "01101010110101111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011000001";
   IN2_i <= "01111000110011000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010111010";
   IN2_i <= "01000100010101010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011101001";
   IN2_i <= "00000101000011011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011011001";
   IN2_i <= "01110100011101001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101100100";
   IN2_i <= "00101100110001110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100010001";
   IN2_i <= "01010110100000011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001010110";
   IN2_i <= "00011100100011111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100110000";
   IN2_i <= "00111010010100110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011010001";
   IN2_i <= "00001111001110101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101010110";
   IN2_i <= "01110001001110010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001001000";
   IN2_i <= "01010011011010101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110001100";
   IN2_i <= "00110101111001010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111000000";
   IN2_i <= "00000110110111101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010110011";
   IN2_i <= "00111001111011011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000001101";
   IN2_i <= "00101101100111000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000111110";
   IN2_i <= "01001110000001110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000010001";
   IN2_i <= "00111100001001001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011111111";
   IN2_i <= "00011111100011101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111000011";
   IN2_i <= "00011011100010110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010010001";
   IN2_i <= "00001110111101010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100010101";
   IN2_i <= "01000110011100110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011011000";
   IN2_i <= "00001000111111101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100000110";
   IN2_i <= "00111101000110001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011001100";
   IN2_i <= "01010111010101101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100100010";
   IN2_i <= "01101000100011001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100010101";
   IN2_i <= "00110011011100001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110111000";
   IN2_i <= "01100110001101000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011001110";
   IN2_i <= "01101001011011101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011011100";
   IN2_i <= "00010000010001111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011011111";
   IN2_i <= "00001111001110001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110000100";
   IN2_i <= "01011010111011010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100101101";
   IN2_i <= "00010000011110001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011000";
   IN2_i <= "00000101110110001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111010011";
   IN2_i <= "00111101001001111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010011110";
   IN2_i <= "00000001001110110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101100011";
   IN2_i <= "00001100000100100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010011111";
   IN2_i <= "01001011001101101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001001110";
   IN2_i <= "01101010000111101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011101000";
   IN2_i <= "01010101001011110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111101111";
   IN2_i <= "01011000110011111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111010111";
   IN2_i <= "00010000110010001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010111";
   IN2_i <= "01100100111011101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010011100";
   IN2_i <= "00101100110111001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010101111";
   IN2_i <= "00100111001111001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111000001";
   IN2_i <= "01101000101001001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001100010";
   IN2_i <= "01001100111101110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111010011";
   IN2_i <= "00110011110010001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000101111";
   IN2_i <= "01001101100110110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011110110";
   IN2_i <= "00100010100100010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000001000";
   IN2_i <= "00111001100011000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110100001";
   IN2_i <= "00111111110000101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010110000";
   IN2_i <= "00100001010000011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010001111";
   IN2_i <= "01100100000100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010110010";
   IN2_i <= "01001001000111001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010100111";
   IN2_i <= "00001101111001101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101111110";
   IN2_i <= "00100010010110001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011000111";
   IN2_i <= "01010011010101101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010101011";
   IN2_i <= "00100101101001001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011100101";
   IN2_i <= "00000110000011111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100101010";
   IN2_i <= "01110100010011000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001000000";
   IN2_i <= "00000001110000101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110000010";
   IN2_i <= "00010111010101111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000110011";
   IN2_i <= "00100101001011110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011011001";
   IN2_i <= "01101000001001011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001111000";
   IN2_i <= "00101101011010010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100101011";
   IN2_i <= "01000001000000001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011000111";
   IN2_i <= "01000011001000100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010001011";
   IN2_i <= "00000010111010111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001011010";
   IN2_i <= "01000010001001011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000110111";
   IN2_i <= "01001000000110010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111001";
   IN2_i <= "01111110001001100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101110000";
   IN2_i <= "01100010010000101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001111010";
   IN2_i <= "00010110011101001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101101110";
   IN2_i <= "01100110101111011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011010001";
   IN2_i <= "01000011010101010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110011111";
   IN2_i <= "00111100111000001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111000100";
   IN2_i <= "01100111001111000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001101101";
   IN2_i <= "01001111110010010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100011011";
   IN2_i <= "01110110101100001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001111";
   IN2_i <= "01111100100101000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011000100";
   IN2_i <= "01101111001111111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100101111";
   IN2_i <= "01101111010000110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010111110";
   IN2_i <= "01110110110110111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110111";
   IN2_i <= "00001010111000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110111010";
   IN2_i <= "00111010111000111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000000101";
   IN2_i <= "01110011000011000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000010001";
   IN2_i <= "01010100000001101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111000000";
   IN2_i <= "00010010010100101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001010011";
   IN2_i <= "00010001000010111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110011001";
   IN2_i <= "01011010011111101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101000010";
   IN2_i <= "01011110101101001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111111011";
   IN2_i <= "00000000110110001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110101111";
   IN2_i <= "00011001010100100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000000100";
   IN2_i <= "01001010101111110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000001100";
   IN2_i <= "00110011000000111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100111011";
   IN2_i <= "01110110101001000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111001111";
   IN2_i <= "00111101111100110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000110101";
   IN2_i <= "00001100100100001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110110011";
   IN2_i <= "01010100011011011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011100011";
   IN2_i <= "01111000011000111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010000000";
   IN2_i <= "01101001001101110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000110000";
   IN2_i <= "00001110000101000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110100001";
   IN2_i <= "01111100111010111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110000";
   IN2_i <= "01000001110110110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100010011";
   IN2_i <= "00001011100101101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111110011";
   IN2_i <= "01100000000001001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100111010";
   IN2_i <= "00101111010000010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000010100";
   IN2_i <= "01100011011110010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011101110";
   IN2_i <= "01111000011111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101101010";
   IN2_i <= "01010010101101100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001001001";
   IN2_i <= "00001001111000110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001011011";
   IN2_i <= "00110100010110011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101011100";
   IN2_i <= "00101010101101010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010011011";
   IN2_i <= "01101001110110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110111101";
   IN2_i <= "00110100110101110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010111111";
   IN2_i <= "01011011101010010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001110011";
   IN2_i <= "01010100001000001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100101010";
   IN2_i <= "00110100001010110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000100100";
   IN2_i <= "00110110010000110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100100100";
   IN2_i <= "00110100010010111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000111100";
   IN2_i <= "01101111101001110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100111001";
   IN2_i <= "01100010010100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011011111";
   IN2_i <= "00000100110011000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001110000";
   IN2_i <= "01101000101101010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111111101";
   IN2_i <= "00100110100111010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010100111";
   IN2_i <= "00100101110100100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010101011";
   IN2_i <= "00100001010110111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110100001";
   IN2_i <= "01110010100110101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010111010";
   IN2_i <= "00110011101000101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010010101";
   IN2_i <= "01001001011010111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100100101";
   IN2_i <= "01011111111100000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001111100";
   IN2_i <= "00111010010010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000001110";
   IN2_i <= "01101001010001001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101100000";
   IN2_i <= "00001100010001001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001000000";
   IN2_i <= "01101110111010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001001101";
   IN2_i <= "01011100011111110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111000000";
   IN2_i <= "01000001001000001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111010001";
   IN2_i <= "00100100110011100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000111011";
   IN2_i <= "00110100111100101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011011010";
   IN2_i <= "01011011100101101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110100010";
   IN2_i <= "01010101100110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101100110";
   IN2_i <= "00001101010110100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111000101";
   IN2_i <= "01010011111001000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000100";
   IN2_i <= "00010100110111011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000111110";
   IN2_i <= "01000001001110010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100111111";
   IN2_i <= "00010011110011111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100010010";
   IN2_i <= "00001110111101010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110100000";
   IN2_i <= "01010010111001100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001001101";
   IN2_i <= "01110110011001111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100111000";
   IN2_i <= "00100001110110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111111100";
   IN2_i <= "00001111110110001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010000111";
   IN2_i <= "00010010011101010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101100110";
   IN2_i <= "01000010101011100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010011000";
   IN2_i <= "00000001011000001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100101101";
   IN2_i <= "01110001010101101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110111001";
   IN2_i <= "01100001101101101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000110";
   IN2_i <= "00001110011101101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010101101";
   IN2_i <= "00011101000010010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101101100";
   IN2_i <= "01000111000100111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001010101";
   IN2_i <= "00001001100010111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010100010";
   IN2_i <= "00111110000010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010011000";
   IN2_i <= "01001001000010100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101001011";
   IN2_i <= "00100101110101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010011";
   IN2_i <= "00111011011000000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001100110";
   IN2_i <= "00100100001001000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011111101";
   IN2_i <= "00111001100111100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100100011";
   IN2_i <= "01110100010111011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010100111";
   IN2_i <= "01111001110101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100100010";
   IN2_i <= "00101010000110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110011111";
   IN2_i <= "01001001000001000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001001100";
   IN2_i <= "00101110001110000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101111101";
   IN2_i <= "01001010110100101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001101111";
   IN2_i <= "00111001101010101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100110101";
   IN2_i <= "00001011011111100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001101";
   IN2_i <= "01110110101111110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100001001";
   IN2_i <= "00000001000101011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000011111";
   IN2_i <= "01010110111110001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101100011";
   IN2_i <= "01001000110100010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000011100";
   IN2_i <= "00110011011100110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101110001";
   IN2_i <= "00110100111111001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010111100";
   IN2_i <= "01011111110110001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101001001";
   IN2_i <= "00001011100010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011101110";
   IN2_i <= "00011111100001000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001011000";
   IN2_i <= "01011100110001000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100110001";
   IN2_i <= "00000000100101110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101010110";
   IN2_i <= "00101100111011001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010101";
   IN2_i <= "01110101111111110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000000000";
   IN2_i <= "00000010011101111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101111101";
   IN2_i <= "01000001010001101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000011001";
   IN2_i <= "01100001001100110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100111010";
   IN2_i <= "00110101110000111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100100010";
   IN2_i <= "01010001110011011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000000";
   IN2_i <= "01100110011011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101101111";
   IN2_i <= "00000010001100011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111110001";
   IN2_i <= "01010011000101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111101110";
   IN2_i <= "01111000110111101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111101100";
   IN2_i <= "01000100110110011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001111111";
   IN2_i <= "01111001101110111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000011000";
   IN2_i <= "01011100110111011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100011";
   IN2_i <= "01101111011001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101100000";
   IN2_i <= "00010111011010000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000000111";
   IN2_i <= "00110101101001101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000111101";
   IN2_i <= "01101111110001100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100010110";
   IN2_i <= "00010101111010101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110011010";
   IN2_i <= "00010000001000000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111011010";
   IN2_i <= "00110001110011101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011100111";
   IN2_i <= "00000100011110101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010011010";
   IN2_i <= "00111101000011011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011111001";
   IN2_i <= "01011011011011111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010111101";
   IN2_i <= "00011110011101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001010011";
   IN2_i <= "00010101010111110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001110101";
   IN2_i <= "01110011001011111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111000001";
   IN2_i <= "00101011111011100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111100";
   IN2_i <= "00101000000000000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010001000";
   IN2_i <= "00000010000111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101010100";
   IN2_i <= "01111110000001001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000000110";
   IN2_i <= "01000010100001010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010000110";
   IN2_i <= "01110010110001101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111000000";
   IN2_i <= "01111001110011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101110000";
   IN2_i <= "00111011000100010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010011001";
   IN2_i <= "00000001010010010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101010111";
   IN2_i <= "00110111000101111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110111010";
   IN2_i <= "00000100010101111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110101100";
   IN2_i <= "00000110000000001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000111011";
   IN2_i <= "00111100110101101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001101000";
   IN2_i <= "00010100100101111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001011010";
   IN2_i <= "01100101111000111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111011111";
   IN2_i <= "01001000000100101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100100100";
   IN2_i <= "01000000001011111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001101010";
   IN2_i <= "01101000111110110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100001000";
   IN2_i <= "00010011010010110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000000111";
   IN2_i <= "01111000101000110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111011001";
   IN2_i <= "01111100000100011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000110000";
   IN2_i <= "00100001010111010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101001001";
   IN2_i <= "00000100100110001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000110001";
   IN2_i <= "01101101010111000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011011111";
   IN2_i <= "01110101001000011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001000101";
   IN2_i <= "01011110100110111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000110001";
   IN2_i <= "00111100011000111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000001010";
   IN2_i <= "00011100110110000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101110";
   IN2_i <= "00101001111100101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010011111";
   IN2_i <= "00010001111010101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001111011";
   IN2_i <= "01101001001001001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111111101";
   IN2_i <= "00010011000011011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110100110";
   IN2_i <= "01011111010001011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010010101";
   IN2_i <= "01001100000110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010010100";
   IN2_i <= "00110001110100010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111000011";
   IN2_i <= "01111010011000111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101100111";
   IN2_i <= "01000111100011010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000010111";
   IN2_i <= "01011111010001101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100010000";
   IN2_i <= "01100001111010100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000011111";
   IN2_i <= "01010111000110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010001111";
   IN2_i <= "00001011111111011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100101111";
   IN2_i <= "01011000110101110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101010001";
   IN2_i <= "00011101001110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111111110";
   IN2_i <= "00100000111011000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001100101";
   IN2_i <= "01011000010101101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001001001";
   IN2_i <= "01011101100101000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110011110";
   IN2_i <= "01010000101101110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010001110";
   IN2_i <= "00100110110101101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100000000";
   IN2_i <= "00001101100011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000001000";
   IN2_i <= "01100011111001001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110000011";
   IN2_i <= "00000100000101110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111110111";
   IN2_i <= "01111011011000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100010111";
   IN2_i <= "01100110101111101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010110100";
   IN2_i <= "01110000111101010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100100001";
   IN2_i <= "00010111011001111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010011";
   IN2_i <= "01100001111000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101101000";
   IN2_i <= "00001001101110011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100111110";
   IN2_i <= "00111100100111011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000001000";
   IN2_i <= "00011010101011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011001000";
   IN2_i <= "00011011110000100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011101";
   IN2_i <= "00101101110001011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000011000";
   IN2_i <= "00110111101100100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101110000";
   IN2_i <= "00011101101001111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010110000";
   IN2_i <= "01010111100110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010001110";
   IN2_i <= "01000000001111011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011010100";
   IN2_i <= "01100000001000111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000010000";
   IN2_i <= "00001111011110000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001111111";
   IN2_i <= "01010101011000110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100010110";
   IN2_i <= "00101011100001101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010000101";
   IN2_i <= "01100110000000011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111001011";
   IN2_i <= "01011101110010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111001011";
   IN2_i <= "00101100100100100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100001111";
   IN2_i <= "01101110111010010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001110";
   IN2_i <= "01100010101011110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010101101";
   IN2_i <= "00010011000010010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011000110";
   IN2_i <= "00001100001011100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100000001";
   IN2_i <= "00011011010100001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100011";
   IN2_i <= "00001111101010101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110111100";
   IN2_i <= "00010010000001000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000010001";
   IN2_i <= "01010111101111011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010111100";
   IN2_i <= "00000011001000000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010111010";
   IN2_i <= "00111011110010011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001010001";
   IN2_i <= "00110001100011110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111101010";
   IN2_i <= "01110110011011100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110110";
   IN2_i <= "00011000011101011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011001101";
   IN2_i <= "00110110110001110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010001010";
   IN2_i <= "01000011010010111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010010010";
   IN2_i <= "01001111101010111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101000110";
   IN2_i <= "00000001111100011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110000";
   IN2_i <= "00100101001101101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110100000";
   IN2_i <= "00000100111110000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001101101";
   IN2_i <= "00111100101010011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010100000";
   IN2_i <= "01110101100011110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101010101";
   IN2_i <= "00101010011100111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010100000";
   IN2_i <= "01010000100010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011110011";
   IN2_i <= "00110110110110110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101101";
   IN2_i <= "00001001010111000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000010110";
   IN2_i <= "00010100101111110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110111010";
   IN2_i <= "00011011100111101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001101110";
   IN2_i <= "00001101110100100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110111";
   IN2_i <= "01001110010001101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101111101";
   IN2_i <= "00110100010111111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010010";
   IN2_i <= "00101010000101011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111000010";
   IN2_i <= "01011100101101011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110011101";
   IN2_i <= "01101001001110101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011101000";
   IN2_i <= "00111100001010001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001100111";
   IN2_i <= "00000000101101100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010101000";
   IN2_i <= "00000011100111010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101100";
   IN2_i <= "01101001110111101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010000101";
   IN2_i <= "00000100010110111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101000000";
   IN2_i <= "00110000100101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101110010";
   IN2_i <= "01100100001001110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010111110";
   IN2_i <= "01011011000011101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000101101";
   IN2_i <= "00111111111011101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011010110";
   IN2_i <= "00110101100011101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001011111";
   IN2_i <= "01111111110010110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000011000";
   IN2_i <= "00011100010101100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111001001";
   IN2_i <= "01001010001010101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000011000";
   IN2_i <= "01010110011111111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001001000";
   IN2_i <= "00111110001101101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011111";
   IN2_i <= "00000111001010000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001110000";
   IN2_i <= "00010000111001011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101010101";
   IN2_i <= "01110011101101111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111000001";
   IN2_i <= "00111011000111001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011000111";
   IN2_i <= "00011011110100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010100111";
   IN2_i <= "00010001000111100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000000000";
   IN2_i <= "01000100101011000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001000";
   IN2_i <= "01010110100110000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110100000";
   IN2_i <= "00101111001000100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011011001";
   IN2_i <= "00111101110100101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011000100";
   IN2_i <= "01001110110110100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100100111";
   IN2_i <= "00101000101011110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000010010";
   IN2_i <= "01001111111101001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100111010";
   IN2_i <= "00010000011001010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111100101";
   IN2_i <= "01100011000111111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000000111";
   IN2_i <= "01000000010100011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110011100";
   IN2_i <= "01001100011011101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000010111";
   IN2_i <= "01000110110010001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000100111";
   IN2_i <= "00101101100100010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000001111";
   IN2_i <= "01010001010001010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000001001";
   IN2_i <= "00110100001100001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000101100";
   IN2_i <= "01011111111010110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001100011";
   IN2_i <= "01000111001001101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011011100";
   IN2_i <= "01010100110110011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111010100";
   IN2_i <= "00010101011001011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001100101";
   IN2_i <= "01110101111100110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011111010";
   IN2_i <= "00110111001011000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011010010";
   IN2_i <= "00000000110110100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000001100";
   IN2_i <= "00111110110101011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000110100";
   IN2_i <= "01101001010111110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011010110";
   IN2_i <= "01000101000100100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010111011";
   IN2_i <= "01101100111110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010011010";
   IN2_i <= "00010011000101011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000100";
   IN2_i <= "01100001011111100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100100111";
   IN2_i <= "01001101001100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001011110";
   IN2_i <= "00101110000001001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000110010";
   IN2_i <= "01100011000001111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010011110";
   IN2_i <= "00111101010000010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110111101";
   IN2_i <= "01101101101010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000000111";
   IN2_i <= "00111011001010100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111100111";
   IN2_i <= "00111011010110110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010111100";
   IN2_i <= "01011100101001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111110111";
   IN2_i <= "01111101001000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000100001";
   IN2_i <= "01001110101001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111001100";
   IN2_i <= "01111100001101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110010010";
   IN2_i <= "01010100110101000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111011";
   IN2_i <= "00111001001000011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110010100";
   IN2_i <= "00101001110011111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011111010";
   IN2_i <= "00001010000101111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001100010";
   IN2_i <= "01000000111000011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100001";
   IN2_i <= "00011010110000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001110100";
   IN2_i <= "00111011000101011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110100010";
   IN2_i <= "01111101010010010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001010110";
   IN2_i <= "01101101001110010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111011000";
   IN2_i <= "01000111110101010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111011110";
   IN2_i <= "01000010110000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011011111";
   IN2_i <= "01110100111110111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101000100";
   IN2_i <= "01010101000100010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011101";
   IN2_i <= "00010011101101111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110111111";
   IN2_i <= "01100110000111110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011001011";
   IN2_i <= "00111010101001110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000100000";
   IN2_i <= "00000100011010111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101001101";
   IN2_i <= "00011110010001110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111100010";
   IN2_i <= "01111001000110100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010011010";
   IN2_i <= "01010000001011100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101110110";
   IN2_i <= "01010101010000100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010000110";
   IN2_i <= "01111101011001110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111110011";
   IN2_i <= "01101011100010001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011000100";
   IN2_i <= "00111001001011110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001010111";
   IN2_i <= "00010100110010010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100001111";
   IN2_i <= "01001101000110000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010001";
   IN2_i <= "01011110001100000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101110";
   IN2_i <= "01011001101000111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000110111";
   IN2_i <= "01111010010111010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000000000";
   IN2_i <= "01001111000010110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010001101";
   IN2_i <= "01011001101111001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100111010";
   IN2_i <= "00101000000100001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111010011";
   IN2_i <= "00101011101110010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000111110";
   IN2_i <= "01110011101000000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110000010";
   IN2_i <= "01000110011101011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000010110";
   IN2_i <= "01101001001011110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100100111";
   IN2_i <= "00101000100000011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011100001";
   IN2_i <= "00110000111010101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101001001";
   IN2_i <= "01000110010001101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101000011";
   IN2_i <= "01111001100110000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101111010";
   IN2_i <= "00111101111111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110010100";
   IN2_i <= "01101101000111110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010101010";
   IN2_i <= "01110011100101100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110000000";
   IN2_i <= "01110001001011011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100000";
   IN2_i <= "00001010000100000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001011101";
   IN2_i <= "00011111011110011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001010101";
   IN2_i <= "00001111111110010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100011100";
   IN2_i <= "01011101010010110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100111101";
   IN2_i <= "00110011101100011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111011011";
   IN2_i <= "01111111000000101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000111011";
   IN2_i <= "00000101110001010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001001110";
   IN2_i <= "01001001001001110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100011001";
   IN2_i <= "01010011010101110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111111110";
   IN2_i <= "00011000010010100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000101010";
   IN2_i <= "00110001001100101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010000010";
   IN2_i <= "01101010110110110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101111001";
   IN2_i <= "01011000110000101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110110001";
   IN2_i <= "01011101111011011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001111110";
   IN2_i <= "01010011000101001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110000101";
   IN2_i <= "01101101001111110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000100001";
   IN2_i <= "01100111000000111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000011101";
   IN2_i <= "01010110001011101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111010111";
   IN2_i <= "00111000010100111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011001001";
   IN2_i <= "01010011110000110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110101111";
   IN2_i <= "01100110010000100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110010";
   IN2_i <= "01010010001110001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110011101";
   IN2_i <= "00000110001010100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000100001";
   IN2_i <= "01110000011111010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010110011";
   IN2_i <= "00011110111110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100101010";
   IN2_i <= "01010000001110000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100010110";
   IN2_i <= "00110010011000001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000011110";
   IN2_i <= "00000011001111111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111000011";
   IN2_i <= "01011110000010000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100110";
   IN2_i <= "00111100101001100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100001100";
   IN2_i <= "00110001100010011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000111011";
   IN2_i <= "01100100001110101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101110110";
   IN2_i <= "01001100110010011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101111011";
   IN2_i <= "00001111001000010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010101000";
   IN2_i <= "01000000001001101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101011010";
   IN2_i <= "01100001001100111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100111";
   IN2_i <= "00011001101110101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001100100";
   IN2_i <= "01000010010111001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110110111";
   IN2_i <= "00011101111010011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011110110";
   IN2_i <= "01001110111001001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111001001";
   IN2_i <= "00001101110010010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101001110";
   IN2_i <= "01101110010110011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010111";
   IN2_i <= "00010010011000010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100001101";
   IN2_i <= "01010100001111000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101100";
   IN2_i <= "01000110111110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010001111";
   IN2_i <= "00110011001000100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100100";
   IN2_i <= "01001000111000110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110100111";
   IN2_i <= "00101110101100001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000111110";
   IN2_i <= "00101010111011010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010011100";
   IN2_i <= "00011101101011001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000110010";
   IN2_i <= "01000111100101001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001010000";
   IN2_i <= "00001110010010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000100110";
   IN2_i <= "00000101001101001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000100011";
   IN2_i <= "00101010100010000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101010001";
   IN2_i <= "00010001011000101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110101000";
   IN2_i <= "00111101001001111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000100";
   IN2_i <= "01001111001000101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000001001";
   IN2_i <= "00111000010101000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010111001";
   IN2_i <= "01000100000001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011111100";
   IN2_i <= "00111011010001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100000110";
   IN2_i <= "01111101010110001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111011101";
   IN2_i <= "01001001000111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101000";
   IN2_i <= "01001100000001101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110011110";
   IN2_i <= "00101011111010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110001000";
   IN2_i <= "00111001111001010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011000110";
   IN2_i <= "00101010011010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000110001";
   IN2_i <= "01000101110111111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110000111";
   IN2_i <= "00000111010011011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011011";
   IN2_i <= "00101111000111001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010001001";
   IN2_i <= "00101000100001100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011110000";
   IN2_i <= "00100111101110100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110011111";
   IN2_i <= "01111011000111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011000011";
   IN2_i <= "01100001110101011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011101110";
   IN2_i <= "01011010001111000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000010011";
   IN2_i <= "00101101011011101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110000001";
   IN2_i <= "01011010111000110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111110010";
   IN2_i <= "00000011001010110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110001110";
   IN2_i <= "01101001101111100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000000011";
   IN2_i <= "01001011110011111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100101011";
   IN2_i <= "01001100010101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110101100";
   IN2_i <= "00000000010101010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001010011";
   IN2_i <= "01010111101101111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111011010";
   IN2_i <= "00001100010101110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100100010";
   IN2_i <= "00100011111000001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100111110";
   IN2_i <= "00001000010101011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101011111";
   IN2_i <= "01100111111100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110100111";
   IN2_i <= "01010101100010011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010000010";
   IN2_i <= "00101101010010000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000010000";
   IN2_i <= "00001010001010101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010101100";
   IN2_i <= "00110100111000000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010101111";
   IN2_i <= "00111011111010001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001000000";
   IN2_i <= "00000101101110010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100100";
   IN2_i <= "00001100010000101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101111001";
   IN2_i <= "01111111010011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000110011";
   IN2_i <= "00011111011111011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000001000";
   IN2_i <= "01010011001101111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110100110";
   IN2_i <= "01111110011001100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101001100";
   IN2_i <= "01011111010100111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110100110";
   IN2_i <= "01011111010001100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001011010";
   IN2_i <= "01110000010001011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100111100";
   IN2_i <= "00110000101010010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100001010";
   IN2_i <= "00001111100110010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010011001";
   IN2_i <= "01110111110110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101010110";
   IN2_i <= "01101010001101101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110101100";
   IN2_i <= "01110100001010010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110111";
   IN2_i <= "01000110011011011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101011101";
   IN2_i <= "00111110010000111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001010010";
   IN2_i <= "01100000111000010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111110101";
   IN2_i <= "01110011101000011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000001101";
   IN2_i <= "01101011000111101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010111001";
   IN2_i <= "00100010100000001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101100011";
   IN2_i <= "01101100110001111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111101110";
   IN2_i <= "00001000001100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010110011";
   IN2_i <= "01111111010101101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011011111";
   IN2_i <= "00110001101100011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001000111";
   IN2_i <= "01001110000111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010100100";
   IN2_i <= "01010100101100010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110110100";
   IN2_i <= "01101010000110101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110111001";
   IN2_i <= "00101110001111010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010001011";
   IN2_i <= "00111000100011100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000010111";
   IN2_i <= "00101001110100110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001101011";
   IN2_i <= "01100001100010111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000111110";
   IN2_i <= "01111000001111000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111100111";
   IN2_i <= "01101110101111111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010011101";
   IN2_i <= "00011110001101111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111101001";
   IN2_i <= "01110101000101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011001100";
   IN2_i <= "01101100100101110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110011110";
   IN2_i <= "00010110100101111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000101011";
   IN2_i <= "00100101100010101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111110100";
   IN2_i <= "00101111100101110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110100001";
   IN2_i <= "01110111001110110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111111000";
   IN2_i <= "00000111000100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000110000";
   IN2_i <= "00000011110010101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110110101";
   IN2_i <= "00000100111011100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101101110";
   IN2_i <= "00000101100110101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101101000";
   IN2_i <= "00110101000100000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100101111";
   IN2_i <= "01000101110110011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101001000";
   IN2_i <= "00101100100100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100110100";
   IN2_i <= "01111111011111000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000011000";
   IN2_i <= "00000011101011001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001110";
   IN2_i <= "01110110000000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000011111";
   IN2_i <= "00100101100000100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110010";
   IN2_i <= "01010100111010000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101101000";
   IN2_i <= "00010100101110111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011000100";
   IN2_i <= "01000100000000110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110011101";
   IN2_i <= "01001010001001101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101001001";
   IN2_i <= "01001101011011001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000110101";
   IN2_i <= "00100001010010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100100100";
   IN2_i <= "01101101000110110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011000110";
   IN2_i <= "00010110010110111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000011011";
   IN2_i <= "00010110011110001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000100010";
   IN2_i <= "01101100111111101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000100000";
   IN2_i <= "00111000000001001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101001101";
   IN2_i <= "01000000110111100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001000010";
   IN2_i <= "00101010100111001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111110001";
   IN2_i <= "01111000110101000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101100010";
   IN2_i <= "01011001011111000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010101100";
   IN2_i <= "00101111101011101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101100100";
   IN2_i <= "01110100100000100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011100000";
   IN2_i <= "00000100111111010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110110011";
   IN2_i <= "01000110001100011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000101110";
   IN2_i <= "01000110010110101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101000000";
   IN2_i <= "01100110100110111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110011001";
   IN2_i <= "00011000011000100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010110000";
   IN2_i <= "00010110110100001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010110111";
   IN2_i <= "00000111001101001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010100000";
   IN2_i <= "00001000010110110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010100101";
   IN2_i <= "00111100010100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110000010";
   IN2_i <= "01100011100101111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100010011";
   IN2_i <= "01011101001100111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110000011";
   IN2_i <= "00101010011001100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110110100";
   IN2_i <= "01001110110101001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111111010";
   IN2_i <= "00011001100110100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010100011";
   IN2_i <= "01110010010000100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011000110";
   IN2_i <= "00010010010111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000001110";
   IN2_i <= "01111100111000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110001100";
   IN2_i <= "00000000011001100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010111000";
   IN2_i <= "01100111110010010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011110111";
   IN2_i <= "01101000111110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111110";
   IN2_i <= "01011001001110001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110110010";
   IN2_i <= "01000000111001101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101110101";
   IN2_i <= "01010110000111100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100100010";
   IN2_i <= "00011001101010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101110100";
   IN2_i <= "00101011000110011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001100100";
   IN2_i <= "01001111010100100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001110000";
   IN2_i <= "00011101101010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110011100";
   IN2_i <= "00001110111001011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111100010";
   IN2_i <= "00000011010000011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101110100";
   IN2_i <= "01110000010110011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100001110";
   IN2_i <= "00100101111100000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000110111";
   IN2_i <= "00010001011111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000011101";
   IN2_i <= "00101111011110111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111110110";
   IN2_i <= "00010010010101101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000111110";
   IN2_i <= "00010110110001001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011000010";
   IN2_i <= "01001111001010111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111110001";
   IN2_i <= "00011101101011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000111011";
   IN2_i <= "00001001001110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010101011";
   IN2_i <= "01010001111000001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101001110";
   IN2_i <= "00010111110011101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001001001";
   IN2_i <= "01010111111010110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010101011";
   IN2_i <= "00101010011000100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010000001";
   IN2_i <= "00000111000110111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010010";
   IN2_i <= "00100010011001101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000001000";
   IN2_i <= "00011111110000000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011101";
   IN2_i <= "00111100011101011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101110101";
   IN2_i <= "01010101000100100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100110100";
   IN2_i <= "00111111101010100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111101011";
   IN2_i <= "00100101110110001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110001000";
   IN2_i <= "00101101111110100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011000110";
   IN2_i <= "00001010000001000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101011111";
   IN2_i <= "01001011010011011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011110011";
   IN2_i <= "00101010110111110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100000001";
   IN2_i <= "01111110000010011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000001111";
   IN2_i <= "00101010110110000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111101100";
   IN2_i <= "01110000110001010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101010011";
   IN2_i <= "00000110101111110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101101101";
   IN2_i <= "01011100101110011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101111";
   IN2_i <= "00111100001111010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101011011";
   IN2_i <= "01111110010100111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010000101";
   IN2_i <= "00000000011011110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001100010";
   IN2_i <= "00100010101100100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001110111";
   IN2_i <= "01000011011111101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010100";
   IN2_i <= "00011001011110000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001011011";
   IN2_i <= "01101001100000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000001100";
   IN2_i <= "01100101011100111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001111000";
   IN2_i <= "00101001010110001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001100111";
   IN2_i <= "00001000111010001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011011000";
   IN2_i <= "01001100110111000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011111010";
   IN2_i <= "00011000001101110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111100001";
   IN2_i <= "00110001001111111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101000100";
   IN2_i <= "01000001010011101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100000110";
   IN2_i <= "00110100010011101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000000000";
   IN2_i <= "00011100011100010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101100111";
   IN2_i <= "01010000101011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001000";
   IN2_i <= "00111100010110101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000100";
   IN2_i <= "01111010111000111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001110110";
   IN2_i <= "01100100011010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111110011";
   IN2_i <= "00100000101110010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100011110";
   IN2_i <= "00100010000010010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000101000";
   IN2_i <= "01010100011001010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101110";
   IN2_i <= "01001011010010110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000000100";
   IN2_i <= "00010010011000100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101001100";
   IN2_i <= "01100111011111110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001000101";
   IN2_i <= "01110010101111111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000101111";
   IN2_i <= "00101011111010101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100110001";
   IN2_i <= "00001011100000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010000100";
   IN2_i <= "01100101010100011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000011100";
   IN2_i <= "00000010111100100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111001";
   IN2_i <= "00001000110100010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010101110";
   IN2_i <= "00100111010110100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001101101";
   IN2_i <= "00011000100101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000111001";
   IN2_i <= "01100111010000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100011011";
   IN2_i <= "01001110011000011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100110111";
   IN2_i <= "01110001100000111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010000001";
   IN2_i <= "01111111111011011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110100111";
   IN2_i <= "01110111110000101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011110010";
   IN2_i <= "00010010101100101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101000110";
   IN2_i <= "00001010110100000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110010100";
   IN2_i <= "01100111001000011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001100000";
   IN2_i <= "01001111000101011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101100100";
   IN2_i <= "01101000111110110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011100101";
   IN2_i <= "00010110110111111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100111010";
   IN2_i <= "01000000011101111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100001110";
   IN2_i <= "00011100111100001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101101100";
   IN2_i <= "01011001000001001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001101";
   IN2_i <= "01011000110000100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110111000";
   IN2_i <= "00110111110110000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011101010";
   IN2_i <= "01000111110000101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000110011";
   IN2_i <= "00110100101111010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011111111";
   IN2_i <= "01000010010110110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111011100";
   IN2_i <= "00000100110011111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100110010";
   IN2_i <= "00001101011000011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001011101";
   IN2_i <= "00101110010100000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100110111";
   IN2_i <= "01110111011011011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000000011";
   IN2_i <= "00101111001100010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110100011";
   IN2_i <= "01000011100100101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001010";
   IN2_i <= "00001111010000011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000000101";
   IN2_i <= "00100101100001000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010011010";
   IN2_i <= "00000011011011000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100110110";
   IN2_i <= "00110101100110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110000110";
   IN2_i <= "01011000110101111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011111101";
   IN2_i <= "01011111011011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110101001";
   IN2_i <= "00010010000100101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000000";
   IN2_i <= "00100111011111011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100001111";
   IN2_i <= "01100001000010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111101001";
   IN2_i <= "01000100110110001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101100";
   IN2_i <= "00101001011111000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111101";
   IN2_i <= "01101100111110101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100000100";
   IN2_i <= "01101011011011011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001111011";
   IN2_i <= "00100011011010011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101010001";
   IN2_i <= "01100100110110101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010010010";
   IN2_i <= "01111010011100100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010110101";
   IN2_i <= "00000011010110010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100111010";
   IN2_i <= "01011111010011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101101110";
   IN2_i <= "00010110000010011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110100010";
   IN2_i <= "00000101101011010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100011101";
   IN2_i <= "00011111100110101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000101010";
   IN2_i <= "01000111011001000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101000111";
   IN2_i <= "01111001001010101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101101010";
   IN2_i <= "00000100001111101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010010111";
   IN2_i <= "01000100101111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001010";
   IN2_i <= "01111110011001101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100110001";
   IN2_i <= "01110011000101011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101000000";
   IN2_i <= "00001001000010110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000001010";
   IN2_i <= "01011100010000101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010010011";
   IN2_i <= "00110110110101011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100101000";
   IN2_i <= "00010111110110001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101010011";
   IN2_i <= "01000001110000000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111001011";
   IN2_i <= "01000011011101101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000111110";
   IN2_i <= "01010110111110100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010010000";
   IN2_i <= "00011100110100110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010100101";
   IN2_i <= "01000111010000000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110111011";
   IN2_i <= "01010010001011100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001111000";
   IN2_i <= "01011010010110011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111000";
   IN2_i <= "01110000100101110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110111010";
   IN2_i <= "01011101110111001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011100111";
   IN2_i <= "01100000000100111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110010011";
   IN2_i <= "00111101110111001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011000000";
   IN2_i <= "00101101111010111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010010001";
   IN2_i <= "01101100100010110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011001101";
   IN2_i <= "01111101000010011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110100000";
   IN2_i <= "01001110010010101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011111111";
   IN2_i <= "01101000001110111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001111110";
   IN2_i <= "01111110010001000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110111010";
   IN2_i <= "00101000010111100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010110011";
   IN2_i <= "01100100100001000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011000";
   IN2_i <= "01100101000001110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111001111";
   IN2_i <= "01011000111010100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100111";
   IN2_i <= "00011111001110010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110011011";
   IN2_i <= "01110110111110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000100010";
   IN2_i <= "01100011001100011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011001101";
   IN2_i <= "01010110101011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110111000";
   IN2_i <= "01001100111110011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100011000";
   IN2_i <= "01110001100001100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011100101";
   IN2_i <= "00010111101010011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010111111";
   IN2_i <= "00011011110110110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101000010";
   IN2_i <= "01001111010010001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111111";
   IN2_i <= "01001101100011010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111100101";
   IN2_i <= "00101001001101000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011110010";
   IN2_i <= "01110101111100011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000111001";
   IN2_i <= "01111100101010011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000010001";
   IN2_i <= "01110000011110001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111011110";
   IN2_i <= "01100011100001010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010101010";
   IN2_i <= "01010110000101011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110010111";
   IN2_i <= "01111011010001000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001100000";
   IN2_i <= "00100000111010110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111001001";
   IN2_i <= "01110011101001100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011101110";
   IN2_i <= "01000000101001110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100010101";
   IN2_i <= "01101001100010001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011111000";
   IN2_i <= "00101010010010100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101111101";
   IN2_i <= "00001001111101101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110010110";
   IN2_i <= "00011010111101000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101111000";
   IN2_i <= "01110101101001011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000010110";
   IN2_i <= "00010111001111100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001010010";
   IN2_i <= "00111000000001011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010010";
   IN2_i <= "01111001111011001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000011011";
   IN2_i <= "01100101001001110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011000000";
   IN2_i <= "00001011111001010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000011010";
   IN2_i <= "00101011010111101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101110100";
   IN2_i <= "00001101110100110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100101000";
   IN2_i <= "01111110001000010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010010011";
   IN2_i <= "00100001101011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101100000";
   IN2_i <= "00000101011111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010010100";
   IN2_i <= "01000111000111000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110110010";
   IN2_i <= "01101101110110011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101110001";
   IN2_i <= "00101101000100101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110011100";
   IN2_i <= "01001100011111111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110111001";
   IN2_i <= "01110101011001110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001011111";
   IN2_i <= "01001100100011101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011011001";
   IN2_i <= "01101001000011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000101";
   IN2_i <= "00010000001100010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010100010";
   IN2_i <= "01000000100111101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000010001";
   IN2_i <= "00111110010110100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111001101";
   IN2_i <= "01110000100101101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110101010";
   IN2_i <= "01101001011101101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001100010";
   IN2_i <= "00101010100001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100001111";
   IN2_i <= "01100000110001111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111010110";
   IN2_i <= "00011100101000110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011100001";
   IN2_i <= "01100011001111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011111000";
   IN2_i <= "00010100010110001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100011011";
   IN2_i <= "01010100111011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111010000";
   IN2_i <= "00100110000010010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001000000";
   IN2_i <= "00010010110010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010110001";
   IN2_i <= "01100100101000010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110000000";
   IN2_i <= "00111010010101001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001011000";
   IN2_i <= "01000001011010001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010111010";
   IN2_i <= "01111011001000011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011110101";
   IN2_i <= "01001100111010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011111001";
   IN2_i <= "01110011001101110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111100101";
   IN2_i <= "01001100100101001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110010101";
   IN2_i <= "00111001010100100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010001";
   IN2_i <= "00111111110001001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000101010";
   IN2_i <= "01110110010110000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000111001";
   IN2_i <= "01101101000001010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101100011";
   IN2_i <= "00111110101001111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011110011";
   IN2_i <= "01000011111111100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111110100";
   IN2_i <= "01001111100110110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010011101";
   IN2_i <= "01010000110101011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011110111";
   IN2_i <= "00010110101010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011001000";
   IN2_i <= "00111000000001010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101001011";
   IN2_i <= "01001101101001100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110011001";
   IN2_i <= "01011000111110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011101";
   IN2_i <= "00000000001110100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001101001";
   IN2_i <= "00111111111110111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000100001";
   IN2_i <= "00010011110010110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010001101";
   IN2_i <= "01000010110000111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011000011";
   IN2_i <= "01000010101010110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001101001";
   IN2_i <= "00111010101111011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101000110";
   IN2_i <= "01100110010110010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101001000";
   IN2_i <= "01100110110110100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000011110";
   IN2_i <= "00011011001001000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011000101";
   IN2_i <= "01000001110011101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001000101";
   IN2_i <= "00001010000010101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011111111";
   IN2_i <= "00001100000111001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111111010";
   IN2_i <= "01101011110110100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110001001";
   IN2_i <= "01111010110110011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000111110";
   IN2_i <= "01011100010001001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001101101";
   IN2_i <= "01101001010011101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001011001";
   IN2_i <= "00010010011001101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000001100";
   IN2_i <= "01110100011101010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001110";
   IN2_i <= "00011110111000001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110000100";
   IN2_i <= "01101110111110100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111010";
   IN2_i <= "01011111001110010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001001100";
   IN2_i <= "01011011010001010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011110";
   IN2_i <= "00111001100011111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110100001";
   IN2_i <= "01101001110010111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000110000";
   IN2_i <= "00111111110011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011101001";
   IN2_i <= "01000111111100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101101011";
   IN2_i <= "00100111110000111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010010011";
   IN2_i <= "00110000111001111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100011010";
   IN2_i <= "01111010010100011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111011010";
   IN2_i <= "00010001101111010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100101010";
   IN2_i <= "01001001101101011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111101111";
   IN2_i <= "00000001001100001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101101101";
   IN2_i <= "01001000010101001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011100001";
   IN2_i <= "00010011100111101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001101000";
   IN2_i <= "00010110110011001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001101101";
   IN2_i <= "01001001000001011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000101111";
   IN2_i <= "00001110110110011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110100010";
   IN2_i <= "00010100001000001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110010100";
   IN2_i <= "00111011101101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101010110";
   IN2_i <= "01000011110011011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111000110";
   IN2_i <= "00011011110101100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110110001";
   IN2_i <= "00010101010001000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110000010";
   IN2_i <= "01011000000001010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001110111";
   IN2_i <= "00001000011001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110111111";
   IN2_i <= "00001111010110010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101110010";
   IN2_i <= "00110010111000001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101011001";
   IN2_i <= "00100000011001001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110010011";
   IN2_i <= "01110011001110010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010001111";
   IN2_i <= "01000100011110001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000110010";
   IN2_i <= "00101101110101010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001111100";
   IN2_i <= "01100010011011101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001110110";
   IN2_i <= "00111011111001101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111111011";
   IN2_i <= "01101011111100001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111001001";
   IN2_i <= "01011010110100000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001111111";
   IN2_i <= "01010010011111111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000100011";
   IN2_i <= "00110011111100001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000001101";
   IN2_i <= "01111011100101010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110011111";
   IN2_i <= "01000110101010101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010010110";
   IN2_i <= "00111111100011110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001000111";
   IN2_i <= "01101001101010100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011111011";
   IN2_i <= "01010011010000101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110100";
   IN2_i <= "01010010100101011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101001011";
   IN2_i <= "01001110111010000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100010000";
   IN2_i <= "01110110110110001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001011111";
   IN2_i <= "00111001010101110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110110110";
   IN2_i <= "00111111011100101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101111111";
   IN2_i <= "00100001100101100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011011100";
   IN2_i <= "00011101001010101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001100101";
   IN2_i <= "00000011101100001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101010";
   IN2_i <= "01101000000000110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010010";
   IN2_i <= "00100110101101111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011101110";
   IN2_i <= "00101101010001011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011100010";
   IN2_i <= "01110011000100011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110011101";
   IN2_i <= "00110110101101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001000110";
   IN2_i <= "00000011000000001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011111110";
   IN2_i <= "01011110010010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100000111";
   IN2_i <= "01000100010100000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100011100";
   IN2_i <= "00110001000100001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111001111";
   IN2_i <= "00101111110010001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000110001";
   IN2_i <= "00100010110110111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100010110";
   IN2_i <= "01010000000110101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010011";
   IN2_i <= "01100110000110101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010000";
   IN2_i <= "00101110110010011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011101101";
   IN2_i <= "00100010111110110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001010010";
   IN2_i <= "00000100000000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101011000";
   IN2_i <= "00010001000111000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110001011";
   IN2_i <= "01001011000100100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001110010";
   IN2_i <= "01100011110010010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010001110";
   IN2_i <= "01010100001011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011000010";
   IN2_i <= "01001101101101011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100001011";
   IN2_i <= "01100011001111000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101100110";
   IN2_i <= "01110011111011011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010011100";
   IN2_i <= "01011011101101111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110000100";
   IN2_i <= "00110000100110001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011000011";
   IN2_i <= "00111101000011001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001000110";
   IN2_i <= "01110111001000001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001000100";
   IN2_i <= "00110100111010000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101110111";
   IN2_i <= "01110101011111100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010010";
   IN2_i <= "00110111001101110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100001110";
   IN2_i <= "01111001111011111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110101011";
   IN2_i <= "00000100110011000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110001";
   IN2_i <= "00010010110001011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011011010";
   IN2_i <= "01001110101000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000001100";
   IN2_i <= "01111111111101110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001111010";
   IN2_i <= "00100000101111011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011000010";
   IN2_i <= "01111011000100011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000001000";
   IN2_i <= "01001100000111011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101010100";
   IN2_i <= "01111011101111001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101010110";
   IN2_i <= "01011011111000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000110101";
   IN2_i <= "00011000100001010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110011";
   IN2_i <= "01111001000001010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110100001";
   IN2_i <= "00111101000110100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001010100";
   IN2_i <= "01101111100110011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110000100";
   IN2_i <= "01011100100110001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100000110";
   IN2_i <= "00001101011011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101111100";
   IN2_i <= "00010001111110000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010000000";
   IN2_i <= "01001011011010010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000010110";
   IN2_i <= "00111010010011100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101000";
   IN2_i <= "01001001111010010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001011100";
   IN2_i <= "00110001010001101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001001010";
   IN2_i <= "00111111111010110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011111001";
   IN2_i <= "01101010111101011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010010101";
   IN2_i <= "00111001101101101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111101";
   IN2_i <= "00110100101011011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100000011";
   IN2_i <= "01000001100101101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111001100";
   IN2_i <= "01100101101011100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001001100";
   IN2_i <= "00001001110001100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000111100";
   IN2_i <= "00111001110100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010110001";
   IN2_i <= "01000111011111101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011111110";
   IN2_i <= "00011000000111110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001100001";
   IN2_i <= "01100100010001010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111011001";
   IN2_i <= "01010010001011010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100100101";
   IN2_i <= "01101010010101011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011010011";
   IN2_i <= "00101000010110110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011011110";
   IN2_i <= "01100101111100011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010111";
   IN2_i <= "01000001110010111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000001000";
   IN2_i <= "00111101100100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111010101";
   IN2_i <= "00000010110001000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000000110";
   IN2_i <= "01101010001001100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000100000";
   IN2_i <= "01111111000010001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110100100";
   IN2_i <= "01010111100100110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010111111";
   IN2_i <= "00010111111101111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000001011";
   IN2_i <= "00110100010111101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000100111";
   IN2_i <= "01001010110001100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011010100";
   IN2_i <= "00000101111010000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110111101";
   IN2_i <= "01111010100101010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000100";
   IN2_i <= "00011011110101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010001111";
   IN2_i <= "00010001111000011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100110011";
   IN2_i <= "01011011110101110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100011011";
   IN2_i <= "00101010100111011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010110111";
   IN2_i <= "00001011001100101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010110110";
   IN2_i <= "00110011101111101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110101011";
   IN2_i <= "01001101011101101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011011011";
   IN2_i <= "01011111001001110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001111";
   IN2_i <= "01110000011100100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100001111";
   IN2_i <= "00101100100100011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100110000";
   IN2_i <= "01000001111010011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101001100";
   IN2_i <= "01011000010110100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000000010";
   IN2_i <= "00000001111001100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001100011";
   IN2_i <= "01000110010010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001110111";
   IN2_i <= "00010010000111010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000100100";
   IN2_i <= "01101111110010010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111101110";
   IN2_i <= "00110101001000000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000001010";
   IN2_i <= "00101011010000101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111110111";
   IN2_i <= "01011110110100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001110101";
   IN2_i <= "00001100110001000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101110000";
   IN2_i <= "01110100010111001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011000110";
   IN2_i <= "01110111100100000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000111100";
   IN2_i <= "01010101001100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011100010";
   IN2_i <= "00100101000000111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100011";
   IN2_i <= "00010010001111011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001000000";
   IN2_i <= "01101100010011101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000101111";
   IN2_i <= "00100001000001001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100100";
   IN2_i <= "01100101111101101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010110110";
   IN2_i <= "00010011100100000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101011111";
   IN2_i <= "01010011000110010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100110";
   IN2_i <= "00000000000010011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000010110";
   IN2_i <= "01001010001010100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101000100";
   IN2_i <= "00011000110010101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111111011";
   IN2_i <= "01100110101001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101001";
   IN2_i <= "01110111111000101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001010";
   IN2_i <= "00100010001010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101111";
   IN2_i <= "00000010100111100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011110100";
   IN2_i <= "01001000010000101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111010011";
   IN2_i <= "01111100111100011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000001111";
   IN2_i <= "01111010011101010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011111000";
   IN2_i <= "01111011010100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111110110";
   IN2_i <= "01001000010000000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101010";
   IN2_i <= "00010101101000011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101111011";
   IN2_i <= "00010110001010010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000010011";
   IN2_i <= "01110110000111001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001011001";
   IN2_i <= "01100010111111100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001011011";
   IN2_i <= "00000100111000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111000000";
   IN2_i <= "00101110000101101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100101110";
   IN2_i <= "00110000111111000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111101000";
   IN2_i <= "01001100011000110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011001001";
   IN2_i <= "01011100110000001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100110";
   IN2_i <= "00010010100011111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011010001";
   IN2_i <= "01000101101110111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101110011";
   IN2_i <= "01001010001011111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101011";
   IN2_i <= "01110000110000011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000010010";
   IN2_i <= "01111000000011010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111001100";
   IN2_i <= "01111100110001010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011101101";
   IN2_i <= "01111111001001011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100001000";
   IN2_i <= "00111100101100011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000111010";
   IN2_i <= "01110010111000010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000101100";
   IN2_i <= "00110110011110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011100110";
   IN2_i <= "01100011000110001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001001101";
   IN2_i <= "00011011100111001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001111101";
   IN2_i <= "01111111010011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100010100";
   IN2_i <= "00101110010011100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010011101";
   IN2_i <= "00110101000100000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110011110";
   IN2_i <= "00111000100100010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110111";
   IN2_i <= "00100001001001111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011010101";
   IN2_i <= "00001010111111001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110100110";
   IN2_i <= "00011010110110001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100011";
   IN2_i <= "01111000101001100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011000101";
   IN2_i <= "01101001011000011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111111011";
   IN2_i <= "01011111111000011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000010100";
   IN2_i <= "01010101100011111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111000110";
   IN2_i <= "00011011111001011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000101101";
   IN2_i <= "01100101110001101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111000100";
   IN2_i <= "01011111001100001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010011100";
   IN2_i <= "01001100111001111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101111111";
   IN2_i <= "00100001011001110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011101";
   IN2_i <= "00001010000010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001110111";
   IN2_i <= "01010010011001000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110110000";
   IN2_i <= "01000011010101011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010000111";
   IN2_i <= "01001000011001101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111011000";
   IN2_i <= "01001100111111001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110110110";
   IN2_i <= "00010000001100011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101101000";
   IN2_i <= "00011010010110100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111000101";
   IN2_i <= "01111110010010001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100101110";
   IN2_i <= "00111110110101010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011111";
   IN2_i <= "01100000000001001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101000100";
   IN2_i <= "00111111010010001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010010001";
   IN2_i <= "01100110000011000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000101110";
   IN2_i <= "01111100010111111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000111011";
   IN2_i <= "00011000011101100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110110110";
   IN2_i <= "00001101010100111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110100110";
   IN2_i <= "00110000100110010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101011110";
   IN2_i <= "01110111110100110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001110000";
   IN2_i <= "01011100011111010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001010000";
   IN2_i <= "01111100010000000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010000100";
   IN2_i <= "01000001110110110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011111111";
   IN2_i <= "01110001101100100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000000001";
   IN2_i <= "00010001111111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100010110";
   IN2_i <= "00000100001110101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101101100";
   IN2_i <= "00000100111000011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001000111";
   IN2_i <= "01100101101010010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111110010";
   IN2_i <= "01100001101111111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101111111";
   IN2_i <= "01011011100101011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010001000";
   IN2_i <= "00111001011111100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010001010";
   IN2_i <= "00101000100010110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000101000";
   IN2_i <= "00111010110101010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100101111";
   IN2_i <= "00000111011101001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000101010";
   IN2_i <= "01110000000110100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001110110";
   IN2_i <= "00000100101100101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000000110";
   IN2_i <= "01110011011110000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111111101";
   IN2_i <= "01000000111100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100000000";
   IN2_i <= "00101011001010111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000100100";
   IN2_i <= "01001110111100010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101111111";
   IN2_i <= "01011101010110000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010100110";
   IN2_i <= "00010101001101001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110000001";
   IN2_i <= "00110110000010110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000101101";
   IN2_i <= "00000000010011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000000101";
   IN2_i <= "00110111000000000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111000";
   IN2_i <= "00100010110001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110111101";
   IN2_i <= "00011110110011101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100001100";
   IN2_i <= "01111000111010100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000011100";
   IN2_i <= "00001111000010110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011111101";
   IN2_i <= "01100000101010110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100110010";
   IN2_i <= "01110101110011010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100000010";
   IN2_i <= "00100101001010111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100111101";
   IN2_i <= "00011011001001100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001001011";
   IN2_i <= "00011010011101101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000010000";
   IN2_i <= "00000011001000111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101111010";
   IN2_i <= "01110011001111111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001101000";
   IN2_i <= "00011100100100000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011101101";
   IN2_i <= "01010001101011100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011000";
   IN2_i <= "01010000001001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001011100";
   IN2_i <= "00111001000100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010111100";
   IN2_i <= "01001000110000010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001011011";
   IN2_i <= "01100010010100111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000010100";
   IN2_i <= "01011000001001110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111110001";
   IN2_i <= "01101111000011001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010100111";
   IN2_i <= "00001001100001101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100111000";
   IN2_i <= "00001110100101101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011101111";
   IN2_i <= "00101110000101100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110101111";
   IN2_i <= "01111110010010110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001100";
   IN2_i <= "01100110011010001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010001011";
   IN2_i <= "01101010111101101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010000010";
   IN2_i <= "00111101110111100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111001011";
   IN2_i <= "00101111100011101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000001001";
   IN2_i <= "00100010011101100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100100001";
   IN2_i <= "01110000001010000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101110111";
   IN2_i <= "01110110110011100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111010000";
   IN2_i <= "01110110011000000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001000010";
   IN2_i <= "00000010100001001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100001110";
   IN2_i <= "00000001010100001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110010011";
   IN2_i <= "00000110000110110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001111111";
   IN2_i <= "00101010101110110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001111111";
   IN2_i <= "01101100010010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011000110";
   IN2_i <= "01101110110110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111101000";
   IN2_i <= "00101111101101001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101011";
   IN2_i <= "01110110000000110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111010";
   IN2_i <= "01110011110001011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000001000";
   IN2_i <= "00011111001111011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001111111";
   IN2_i <= "01100011010110011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110111101";
   IN2_i <= "01011010111011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100110011";
   IN2_i <= "00011111100101111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110001110";
   IN2_i <= "00011011101110011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000001011";
   IN2_i <= "00100110100100001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100011010";
   IN2_i <= "00001010010111011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011111011";
   IN2_i <= "00001100111110010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100100101";
   IN2_i <= "01110101010010100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000010";
   IN2_i <= "01101001000101100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110111110";
   IN2_i <= "01101001110101111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000100";
   IN2_i <= "01011111101101010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110110110";
   IN2_i <= "01110101000111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110110100";
   IN2_i <= "00100100011000101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000001011";
   IN2_i <= "00111100110001010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111000101";
   IN2_i <= "00100001010100000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100000111";
   IN2_i <= "01010010011011010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001010001";
   IN2_i <= "01011101000100011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011110000";
   IN2_i <= "00111110000010011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000000001";
   IN2_i <= "00001010000110100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010101101";
   IN2_i <= "01000011111010010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010010000";
   IN2_i <= "00001010111001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101001";
   IN2_i <= "01101111011100011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010100011";
   IN2_i <= "01100000111000110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101011101";
   IN2_i <= "01000101101100001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110011101";
   IN2_i <= "00011100000010101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000110001";
   IN2_i <= "00111011101111000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000001";
   IN2_i <= "01111010010000011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010011010";
   IN2_i <= "00001111010101100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001011";
   IN2_i <= "00101001001000111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100010000";
   IN2_i <= "00001000000001101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101101010";
   IN2_i <= "01110010101011110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110001000";
   IN2_i <= "00100110100010011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101001001";
   IN2_i <= "01101110001101100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100010011";
   IN2_i <= "00001000010111001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110000010";
   IN2_i <= "00101000010111001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111110100";
   IN2_i <= "01110000010011101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000011010";
   IN2_i <= "00110011011111111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111011111";
   IN2_i <= "00010000000101101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101000110";
   IN2_i <= "00001111111001010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011110011";
   IN2_i <= "00101011101110011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001010101";
   IN2_i <= "00111001010111110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110110000";
   IN2_i <= "00010110100100111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000010000";
   IN2_i <= "01010010010010000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101111100";
   IN2_i <= "01001110010111110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010001111";
   IN2_i <= "00011011110110110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111111111";
   IN2_i <= "01000010100101011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110011011";
   IN2_i <= "00101010010010010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101101";
   IN2_i <= "00111010001100001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010010110";
   IN2_i <= "00010111010111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001111001";
   IN2_i <= "00011011111001101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000011001";
   IN2_i <= "01100001001000011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110000100";
   IN2_i <= "01101110000010101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000011110";
   IN2_i <= "01100101111110000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100100";
   IN2_i <= "00000100111110100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101010111";
   IN2_i <= "00111111000010100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101000001";
   IN2_i <= "00100110110001000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000000001";
   IN2_i <= "01100101010110101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110110011";
   IN2_i <= "00010101100100011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011000110";
   IN2_i <= "01000001110011110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111010111";
   IN2_i <= "01111101010011011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110011000";
   IN2_i <= "00001011111110110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101001100";
   IN2_i <= "01101011000101100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100000011";
   IN2_i <= "01111111100111001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011001101";
   IN2_i <= "01001000000101100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000100011";
   IN2_i <= "01001010111101001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101110";
   IN2_i <= "00001100101000000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010100011";
   IN2_i <= "01000000001101100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110000101";
   IN2_i <= "00111110111000100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001001100";
   IN2_i <= "00101011001110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010011110";
   IN2_i <= "01101110100101100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110110010";
   IN2_i <= "01010011000001000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101111110";
   IN2_i <= "01100101110111001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010010001";
   IN2_i <= "01101000011110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100101011";
   IN2_i <= "01001110101001110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110000";
   IN2_i <= "01110011010101110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111101000";
   IN2_i <= "00011101100001000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000111001";
   IN2_i <= "00111110101000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110111";
   IN2_i <= "00110110111001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000001001";
   IN2_i <= "00100110100101001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000001";
   IN2_i <= "01101101111011101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100110";
   IN2_i <= "00110010110011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111100011";
   IN2_i <= "01011101001101110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001010010";
   IN2_i <= "00110000111100101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110101011";
   IN2_i <= "00110001011010111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111011110";
   IN2_i <= "01001000110000010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100111";
   IN2_i <= "00111000110111101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011011111";
   IN2_i <= "00000001000100110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000111111";
   IN2_i <= "01011001110111010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100001111";
   IN2_i <= "00011000001001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100000001";
   IN2_i <= "01101000100110000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101010000";
   IN2_i <= "01100111101010111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010011110";
   IN2_i <= "01001111100011110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011001000";
   IN2_i <= "01110110111110100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110111110";
   IN2_i <= "00011100000110011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011110110";
   IN2_i <= "01001000010011110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111100100";
   IN2_i <= "01100100010000111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101110011";
   IN2_i <= "01111010100111110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001011000";
   IN2_i <= "01100000111001100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000010010";
   IN2_i <= "01101100101100000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111001111";
   IN2_i <= "00110010101011110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111011101";
   IN2_i <= "00100001111010010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011110100";
   IN2_i <= "01100011111100100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111100001";
   IN2_i <= "00100011000010111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010010111";
   IN2_i <= "01110010000101001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010110110";
   IN2_i <= "01101100001001011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100000001";
   IN2_i <= "00110010111000110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101101000";
   IN2_i <= "00101011100110010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101100010";
   IN2_i <= "01010001011011010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110110010";
   IN2_i <= "00111101010100001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110100110";
   IN2_i <= "00000000010011010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110111101";
   IN2_i <= "01011111111010010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111001111";
   IN2_i <= "00100110000000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010111";
   IN2_i <= "00000001000010001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111011111";
   IN2_i <= "00011000110000101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110000001";
   IN2_i <= "00011100111101111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111110000";
   IN2_i <= "01100110111011001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110111010";
   IN2_i <= "00010001000011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010000101";
   IN2_i <= "01111010111000110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100101010";
   IN2_i <= "01011111100101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010110101";
   IN2_i <= "00000000010101011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000111011";
   IN2_i <= "01011000110100011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101010110";
   IN2_i <= "01001011000111100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000111100";
   IN2_i <= "01001010010101010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110111110";
   IN2_i <= "01011000110111000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001111110";
   IN2_i <= "01111101000111000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001001101";
   IN2_i <= "00101000100100011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110011010";
   IN2_i <= "01100001101011111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110011";
   IN2_i <= "00000000101111011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111101110";
   IN2_i <= "00100110110111010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111000100";
   IN2_i <= "01000100111101000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110001110";
   IN2_i <= "01101000101000100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110100100";
   IN2_i <= "01000000000000100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000010001";
   IN2_i <= "01100111110001110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010000100";
   IN2_i <= "01001011110101011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110100011";
   IN2_i <= "01111110110011111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111001011";
   IN2_i <= "00110011111101111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011101110";
   IN2_i <= "01111000101100011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110110110";
   IN2_i <= "01101001011011101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000011110";
   IN2_i <= "00101110111010101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010101011";
   IN2_i <= "00010110110110000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100011111";
   IN2_i <= "01000010011011000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101011111";
   IN2_i <= "01000011101101000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100001";
   IN2_i <= "00110010100010001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010001110";
   IN2_i <= "00100000101100100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110100111";
   IN2_i <= "00000000101100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001111001";
   IN2_i <= "01011010010011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000011101";
   IN2_i <= "01111111110111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110111001";
   IN2_i <= "00110011010111001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110111000";
   IN2_i <= "01011111011011011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101101000";
   IN2_i <= "00110101110101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000000";
   IN2_i <= "01000110010100111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110011110";
   IN2_i <= "00101011100010111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110111111";
   IN2_i <= "00001011111101101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110000111";
   IN2_i <= "00000010000010101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011100";
   IN2_i <= "01100001101110110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011100110";
   IN2_i <= "00011000000101110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011101101";
   IN2_i <= "01101101111101000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111001010";
   IN2_i <= "00011011100100110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110111000";
   IN2_i <= "00110000010011010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111000111";
   IN2_i <= "00100101011100100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110111001";
   IN2_i <= "01011100101010011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011101011";
   IN2_i <= "00011111110110010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110010001";
   IN2_i <= "00000000011001000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001110101";
   IN2_i <= "00100101100010000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000000000";
   IN2_i <= "01010111110000111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010001100";
   IN2_i <= "01001100101011100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010111000";
   IN2_i <= "01010010000010101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011001000";
   IN2_i <= "01110100110011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011100101";
   IN2_i <= "01100100000001101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010111000";
   IN2_i <= "01010110011000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110011001";
   IN2_i <= "00010001111010110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100101001";
   IN2_i <= "00110010001100100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001110000";
   IN2_i <= "00010110011001000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100001";
   IN2_i <= "00111000110010101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101100110";
   IN2_i <= "01000100000101100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100101100";
   IN2_i <= "00110001010011000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000001111";
   IN2_i <= "00001011111101101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101110001";
   IN2_i <= "01111001101010111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100000111";
   IN2_i <= "00100110011011010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111010101";
   IN2_i <= "01011011110011011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011100010";
   IN2_i <= "00101100010001100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100011011";
   IN2_i <= "01111110010001111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010110111";
   IN2_i <= "00100011010101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101111101";
   IN2_i <= "00111010101001011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101100000";
   IN2_i <= "00011011110000010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111101101";
   IN2_i <= "00101110011010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000101";
   IN2_i <= "01101010101010010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010111100";
   IN2_i <= "01101101001101011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001100001";
   IN2_i <= "00111010010111101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100000110";
   IN2_i <= "00100000001110010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011000";
   IN2_i <= "00100000010101100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100001000";
   IN2_i <= "01111111010010111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101111100";
   IN2_i <= "01100000111110010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000111";
   IN2_i <= "01101110001100100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000101101";
   IN2_i <= "01011011001100101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100111000";
   IN2_i <= "00100001011101011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001000100";
   IN2_i <= "01011101111011111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111100100";
   IN2_i <= "00000010011100001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010100110";
   IN2_i <= "01100011100110100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000111111";
   IN2_i <= "01101000010101111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100101";
   IN2_i <= "01101001110010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111110111";
   IN2_i <= "01010110111001110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011100";
   IN2_i <= "00001011011111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010110010";
   IN2_i <= "01111011111101101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111011";
   IN2_i <= "00001101000101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000110001";
   IN2_i <= "00101000011110010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100000100";
   IN2_i <= "01111100111100111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100110000";
   IN2_i <= "01110011001001000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001111000";
   IN2_i <= "00010010010001101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101001100";
   IN2_i <= "01010011010000011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101111100";
   IN2_i <= "01001010101110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010101111";
   IN2_i <= "01011000111010101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011110111";
   IN2_i <= "00110010111111101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111111";
   IN2_i <= "01011000110011001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101010001";
   IN2_i <= "00110101001010100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111010000";
   IN2_i <= "01111011100010100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101100011";
   IN2_i <= "01010001110111010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101011101";
   IN2_i <= "00000110000100100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011001101";
   IN2_i <= "00101010100110010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001110101";
   IN2_i <= "00110011001101000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010111001";
   IN2_i <= "00001001100011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010100101";
   IN2_i <= "00110111101100010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111011111";
   IN2_i <= "01100000111100010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011010100";
   IN2_i <= "00010010000101000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110001101";
   IN2_i <= "00000011111101000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101010110";
   IN2_i <= "00000100010100110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011100110";
   IN2_i <= "00011101001100110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011000011";
   IN2_i <= "00000110100001110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010000011";
   IN2_i <= "00101000101111011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111011";
   IN2_i <= "01100101000100000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001010010";
   IN2_i <= "00001011110001101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101110010";
   IN2_i <= "00110001011111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100011001";
   IN2_i <= "00110011101101011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101101001";
   IN2_i <= "01010000100111110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110101010";
   IN2_i <= "00100001011100111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110110000";
   IN2_i <= "00000010000000010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101100100";
   IN2_i <= "01100100111000100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010011010";
   IN2_i <= "01100110110010001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010000101";
   IN2_i <= "00010110011100110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000101100";
   IN2_i <= "00101011111100011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111010";
   IN2_i <= "00110010101110111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010101010";
   IN2_i <= "00001010110000100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101010";
   IN2_i <= "00101000000100101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001111011";
   IN2_i <= "00111111100110110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000110111";
   IN2_i <= "00100000010100011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001011101";
   IN2_i <= "00001100101000110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001100000";
   IN2_i <= "01000111110011000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000101111";
   IN2_i <= "00100000001110001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111000011";
   IN2_i <= "00111101110000001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000000011";
   IN2_i <= "01111101001000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101001010";
   IN2_i <= "01110011101010100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110101";
   IN2_i <= "01110111110110111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101100000";
   IN2_i <= "01110111111001011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001111111";
   IN2_i <= "01101111001100001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111100010";
   IN2_i <= "01100111000110000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111111100";
   IN2_i <= "01001000000001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100100100";
   IN2_i <= "01000000110011110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100101100";
   IN2_i <= "00000011101100000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101110110";
   IN2_i <= "00011111010000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110100111";
   IN2_i <= "01001001001010000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101101000";
   IN2_i <= "01100111011110011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100101";
   IN2_i <= "00001100001111110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111001111";
   IN2_i <= "01000000000011000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100111";
   IN2_i <= "01100000001011110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101000111";
   IN2_i <= "00011101011111010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000001101";
   IN2_i <= "01001001000111101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110110010";
   IN2_i <= "01010100101000101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101111111";
   IN2_i <= "01101010000111001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101000011";
   IN2_i <= "00001100000110100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010110101";
   IN2_i <= "01000010011110001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111001111";
   IN2_i <= "00011011100110101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101011101";
   IN2_i <= "01010001010001110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011010011";
   IN2_i <= "01111101000010100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100000011";
   IN2_i <= "01011010111100000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101110111";
   IN2_i <= "00101111011010010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110011";
   IN2_i <= "01001100111000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001011001";
   IN2_i <= "00011101110101000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111100010";
   IN2_i <= "00011010000011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111010110";
   IN2_i <= "01101111001100100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100101010";
   IN2_i <= "00100111111110111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101011001";
   IN2_i <= "01101011111110010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010111001";
   IN2_i <= "00110110010001000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110010110";
   IN2_i <= "00101000100011010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010001011";
   IN2_i <= "00110011001110111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000001010";
   IN2_i <= "01111001111011011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010010100";
   IN2_i <= "00000010011010010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101110000";
   IN2_i <= "00111010000110000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011000011";
   IN2_i <= "01000101000001000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111110000";
   IN2_i <= "00001110000010101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000000011";
   IN2_i <= "00101101000100110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101010010";
   IN2_i <= "01111111000001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101010110";
   IN2_i <= "00110110110011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001010011";
   IN2_i <= "00010011010000110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100010111";
   IN2_i <= "01111000101110011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111011101";
   IN2_i <= "01000111110001011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000110010";
   IN2_i <= "00100000101011001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001000001";
   IN2_i <= "01011110100011100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011111000";
   IN2_i <= "01000001101011110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110100001";
   IN2_i <= "00000010001001111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111000111";
   IN2_i <= "01000000011011011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110111111";
   IN2_i <= "01000111111100100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100101111";
   IN2_i <= "01101100100101101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100010101";
   IN2_i <= "01011101100011000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111111110";
   IN2_i <= "01100011110000111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011101000";
   IN2_i <= "01010101001011011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000101101";
   IN2_i <= "01001110011111101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111011110";
   IN2_i <= "01100010001100011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110101101";
   IN2_i <= "00100100110111010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110111010";
   IN2_i <= "01100001101001110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111111001";
   IN2_i <= "00100010011101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010010001";
   IN2_i <= "01010000100111101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111011000";
   IN2_i <= "01110111001111101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001001011";
   IN2_i <= "01001011101100100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101001111";
   IN2_i <= "00100011011010000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101110100";
   IN2_i <= "00100010110011110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100110001";
   IN2_i <= "00111100111101001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101101011";
   IN2_i <= "01110010000110001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000100";
   IN2_i <= "00111001100110101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000010111";
   IN2_i <= "00111110101001000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000010101";
   IN2_i <= "00110100010100001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101111001";
   IN2_i <= "00110011101100111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110011111";
   IN2_i <= "01111101001100000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111000010";
   IN2_i <= "00001110110011111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101000111";
   IN2_i <= "00000110110110110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101001100";
   IN2_i <= "01111101100100000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100111111";
   IN2_i <= "00111001001000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101100011";
   IN2_i <= "00100111000100010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100101010";
   IN2_i <= "01110111101110111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001011000";
   IN2_i <= "01100000101001100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001010010";
   IN2_i <= "01100110010100100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101100010";
   IN2_i <= "00110001010010111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100000011";
   IN2_i <= "01111110011000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011011100";
   IN2_i <= "01110110101110100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100010001";
   IN2_i <= "01100111000111010";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000001110";
   IN2_i <= "01110000001010001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100001010";
   IN2_i <= "01011100110001011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010101010";
   IN2_i <= "01100101000010000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010101101";
   IN2_i <= "01100010011000001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010100011";
   IN2_i <= "00010100011100101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001010011";
   IN2_i <= "01001101000111111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110011000";
   IN2_i <= "01111001001111010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001000100";
   IN2_i <= "00101100001001000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110011101";
   IN2_i <= "00000010001011011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000100100";
   IN2_i <= "00100011011111001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010100010";
   IN2_i <= "00010100011101000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000001010";
   IN2_i <= "01000001110001011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111100011";
   IN2_i <= "00110100100110101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111001110";
   IN2_i <= "00001000000111110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111001";
   IN2_i <= "00101110110111100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110010101";
   IN2_i <= "00001010101100111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111110111";
   IN2_i <= "01110111101110000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111111000";
   IN2_i <= "01001000101101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000010110";
   IN2_i <= "01000011001101010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011100010";
   IN2_i <= "00001111111011110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010011010";
   IN2_i <= "01100100011011100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101101101";
   IN2_i <= "01001111000011001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111010011";
   IN2_i <= "00010011011011001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100000111";
   IN2_i <= "01011011000010010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110100101";
   IN2_i <= "00110000111101100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100001111";
   IN2_i <= "01100100110010100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011010001";
   IN2_i <= "01110010111000010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111001010";
   IN2_i <= "00000111001100110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100110110";
   IN2_i <= "01100011001101111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011100000";
   IN2_i <= "01100111101010111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110101100";
   IN2_i <= "01101010101000111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000111100";
   IN2_i <= "00100100001001110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010111000";
   IN2_i <= "00000011110101100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011010101";
   IN2_i <= "00100001000111111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110101111";
   IN2_i <= "00100101100001101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011111111";
   IN2_i <= "00111000101100101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100111000";
   IN2_i <= "00001001001001011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000010011";
   IN2_i <= "00011010101110101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010000101";
   IN2_i <= "01010110011010000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001110100";
   IN2_i <= "00011110101011010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011110110";
   IN2_i <= "01101000000000111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000101011";
   IN2_i <= "00000001110011010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100110011";
   IN2_i <= "00100101101100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110011110";
   IN2_i <= "01110000001101011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100101110";
   IN2_i <= "00001011000100111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101001111";
   IN2_i <= "00100001101010101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111101011";
   IN2_i <= "01011000000111110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010100111";
   IN2_i <= "00111100011110001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100000111";
   IN2_i <= "00010010100011101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101111011";
   IN2_i <= "00101000010111100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110010100";
   IN2_i <= "01101100101111010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001000110";
   IN2_i <= "00011110110010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110010000";
   IN2_i <= "00100110110001110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111101000";
   IN2_i <= "00101110000011000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101110111";
   IN2_i <= "00100110001100110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001010100";
   IN2_i <= "00111011110100111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000100011";
   IN2_i <= "00111100100111101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101110000";
   IN2_i <= "00100110110000001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001001000";
   IN2_i <= "01100111111110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111111100";
   IN2_i <= "00000011100010111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110111110";
   IN2_i <= "00001010100011100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110011001";
   IN2_i <= "01001001010000100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110101110";
   IN2_i <= "01101111110010001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111111001";
   IN2_i <= "01001010100010011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100111100";
   IN2_i <= "01100111101011111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000100000";
   IN2_i <= "00100010101001000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001000110";
   IN2_i <= "00000010101001001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001001110";
   IN2_i <= "00010011110011110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101111000";
   IN2_i <= "01000010000011010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001000110";
   IN2_i <= "00111010011010010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000110010";
   IN2_i <= "00101111111011011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101111111";
   IN2_i <= "00001011111101101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010100100";
   IN2_i <= "00101111110001000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011100";
   IN2_i <= "01101110100110000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110010000";
   IN2_i <= "00010001010110110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000011010";
   IN2_i <= "00101010110101111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100000000";
   IN2_i <= "01100011110001010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100111100";
   IN2_i <= "01111100001000110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100011101";
   IN2_i <= "01111000001111011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000111110";
   IN2_i <= "01100111101011100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000000111";
   IN2_i <= "00100000010000111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111100111";
   IN2_i <= "01110110000000001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111010111";
   IN2_i <= "01100000001011011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110001100";
   IN2_i <= "00110010010001111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101100110";
   IN2_i <= "01011011010010100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000011010";
   IN2_i <= "00010110011000100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111100111";
   IN2_i <= "00100100101010110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010010011";
   IN2_i <= "00001110110001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001011101";
   IN2_i <= "01000110011000110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110011011";
   IN2_i <= "00101110100100000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101010000";
   IN2_i <= "01100110101011001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110010101";
   IN2_i <= "01001101011111110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011000110";
   IN2_i <= "01101100101111001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000100000";
   IN2_i <= "00010000000110111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100111111";
   IN2_i <= "00011011111101000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010101";
   IN2_i <= "01000010011011011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110101110";
   IN2_i <= "01111111011010010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010000";
   IN2_i <= "00010101011011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100110001";
   IN2_i <= "01010111000100000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011100001";
   IN2_i <= "00101100011001010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111011011";
   IN2_i <= "01010101010011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000111";
   IN2_i <= "00000010000100110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111110000";
   IN2_i <= "00100001001011001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100100011";
   IN2_i <= "00011011111001000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011011000";
   IN2_i <= "00100010000011111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111010111";
   IN2_i <= "00001100111011101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001001010";
   IN2_i <= "01010000001111111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110011000";
   IN2_i <= "01100100111101000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100011";
   IN2_i <= "00111111101100011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101000111";
   IN2_i <= "01101001110100101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000011011";
   IN2_i <= "01100011111101001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100110101";
   IN2_i <= "00000011011101010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001111101";
   IN2_i <= "00111111100011101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100011001";
   IN2_i <= "01011100001011110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010110110";
   IN2_i <= "01010001010100111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101011101";
   IN2_i <= "01100010111001101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011010011";
   IN2_i <= "01111001101111111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001111001";
   IN2_i <= "00101001010010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001101110";
   IN2_i <= "00111110100011011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111011";
   IN2_i <= "01100111111101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000010";
   IN2_i <= "01000100000110000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011001010";
   IN2_i <= "00010100000100111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111100111";
   IN2_i <= "01001010010011000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110001100";
   IN2_i <= "01101100100110101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011010001";
   IN2_i <= "01010001001001010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010000000";
   IN2_i <= "00010000111001110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100011001";
   IN2_i <= "00001100001111010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110011001";
   IN2_i <= "01010110100011001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111111010";
   IN2_i <= "01101110000010010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110010011";
   IN2_i <= "01001101110000100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001000100";
   IN2_i <= "01010001011001010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111011110";
   IN2_i <= "01000000111010100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001111101";
   IN2_i <= "00100110011111111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010111001";
   IN2_i <= "01100101110101000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111010101";
   IN2_i <= "00001001011101101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100000110";
   IN2_i <= "00010110101100111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101000110";
   IN2_i <= "00111110011010000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110101000";
   IN2_i <= "00100011100101010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000111011";
   IN2_i <= "01011101101011110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010010101";
   IN2_i <= "00000110111111100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000111000";
   IN2_i <= "00110001010001010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101110";
   IN2_i <= "00001110100110101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100101010";
   IN2_i <= "00011011111101101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110100";
   IN2_i <= "00111011001110001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001111010";
   IN2_i <= "00000001011111100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101001011";
   IN2_i <= "00100011001011111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101100111";
   IN2_i <= "01001110000111010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011000111";
   IN2_i <= "01101101000010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100000001";
   IN2_i <= "01000011000100101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100101000";
   IN2_i <= "00111101111100101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011000111";
   IN2_i <= "00001101110100101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010111110";
   IN2_i <= "00010111110011111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010000110";
   IN2_i <= "01110111111101101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111011000";
   IN2_i <= "01101000110010001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100010100";
   IN2_i <= "01011100011001000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010111110";
   IN2_i <= "01001000011100011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010110100";
   IN2_i <= "00110001101011110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000110";
   IN2_i <= "00011010000110011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010100111";
   IN2_i <= "01111001110010111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111010011";
   IN2_i <= "01010101000010110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111011";
   IN2_i <= "00111010110011001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001001101";
   IN2_i <= "01111110110010000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100001010";
   IN2_i <= "01100101000011100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111011010";
   IN2_i <= "00010110110111011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011000011";
   IN2_i <= "00101011111010111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110111100";
   IN2_i <= "01011110000011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110011010110";
   IN2_i <= "01011101011101100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001111001";
   IN2_i <= "00001111000001101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111011101";
   IN2_i <= "00011011011000110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100011";
   IN2_i <= "01100101100001001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111100111";
   IN2_i <= "01010001100011001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010000001";
   IN2_i <= "01000000110100100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100101010";
   IN2_i <= "00000010000101000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010011011";
   IN2_i <= "00000111110110111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101101100";
   IN2_i <= "00100001011101101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010100110";
   IN2_i <= "01101010011010111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100011100";
   IN2_i <= "00000001001100000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110111111";
   IN2_i <= "00011010101001100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101101101";
   IN2_i <= "00110001010111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001100011";
   IN2_i <= "01100100010001110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011110010";
   IN2_i <= "00010000111000000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001010010";
   IN2_i <= "00101111001111001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011011000";
   IN2_i <= "01000110100101010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001110001";
   IN2_i <= "00101011001000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111111110";
   IN2_i <= "00101111111100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111101111";
   IN2_i <= "01100010000100111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001100011";
   IN2_i <= "00111000001011110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010000010";
   IN2_i <= "00010001001000110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001111101";
   IN2_i <= "00100001010000110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100001101";
   IN2_i <= "00110000110011001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101001100";
   IN2_i <= "00100110000101011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001000110";
   IN2_i <= "00011010010001110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000111010";
   IN2_i <= "01111111110001010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101110101";
   IN2_i <= "01110110100010110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000111110";
   IN2_i <= "01111111110011000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001000110";
   IN2_i <= "01110011011001010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001110110";
   IN2_i <= "00001100000001000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111010011";
   IN2_i <= "01010101110100000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111101100";
   IN2_i <= "00010001101100101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010001001";
   IN2_i <= "00011101000111100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111110000";
   IN2_i <= "01000001111011000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101011011";
   IN2_i <= "00110111111111000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111010011";
   IN2_i <= "01100011111001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100101100";
   IN2_i <= "01010110111011111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100111000";
   IN2_i <= "00000000000101011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000110110";
   IN2_i <= "00100110011101101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000011110";
   IN2_i <= "00111110100001111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011111";
   IN2_i <= "01010001111110110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111011000";
   IN2_i <= "01010111001011011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111110111";
   IN2_i <= "00111001101101110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110111110";
   IN2_i <= "00110001100010000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000101000";
   IN2_i <= "01001110000000001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011110111";
   IN2_i <= "01101111011001011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101100100";
   IN2_i <= "01100100011101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010110111";
   IN2_i <= "01001101010101111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110010111";
   IN2_i <= "01111001110000100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101010010";
   IN2_i <= "01100110001001011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001010";
   IN2_i <= "00111100000100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111010010";
   IN2_i <= "01100011110000101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010010111";
   IN2_i <= "01001001001010101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110000";
   IN2_i <= "00010110001111001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110000110";
   IN2_i <= "01110101101110011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100101111";
   IN2_i <= "01100001110001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101100";
   IN2_i <= "01000100110110001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011011001";
   IN2_i <= "00000111100100100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010000101";
   IN2_i <= "01011011001101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101010011";
   IN2_i <= "00011110011010000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101001";
   IN2_i <= "01011100011101101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101001000";
   IN2_i <= "01111001110111111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011000000";
   IN2_i <= "00101100011000101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000110100";
   IN2_i <= "00010101011100101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011011010";
   IN2_i <= "01010101101010011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111100";
   IN2_i <= "00101010111110000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111001000";
   IN2_i <= "01110101001111000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111001010";
   IN2_i <= "00000110000000111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110010001";
   IN2_i <= "01100110010110010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010111111";
   IN2_i <= "00101100111001110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010111111";
   IN2_i <= "00000100110000000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100010111";
   IN2_i <= "00001111000110111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000000101";
   IN2_i <= "01101110111010000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001010100";
   IN2_i <= "00111001111111011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000010000";
   IN2_i <= "01000111001110010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110101100";
   IN2_i <= "00101100100001111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111111000";
   IN2_i <= "01001000101101100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100000010";
   IN2_i <= "00010001000000110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100101101";
   IN2_i <= "01011111101011001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100101110";
   IN2_i <= "00100111111100111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001010111";
   IN2_i <= "01101110000101000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010110011";
   IN2_i <= "01001101101010110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111000111";
   IN2_i <= "01010100000110110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001110000";
   IN2_i <= "01110100001111100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010001111";
   IN2_i <= "00001001000010010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010110111";
   IN2_i <= "01110111011010010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101010000";
   IN2_i <= "01011010100001001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001111011";
   IN2_i <= "00000010010101110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001111100";
   IN2_i <= "01001001110010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010101100";
   IN2_i <= "00100101010110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001100100";
   IN2_i <= "01110100110011011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101110101";
   IN2_i <= "00100000000101100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001101110";
   IN2_i <= "01011010100000101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101011111";
   IN2_i <= "01010010111011111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001000000";
   IN2_i <= "01100110100100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101010011";
   IN2_i <= "01011011000001100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001000010";
   IN2_i <= "00101000001110011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001110001";
   IN2_i <= "01001100111001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001011";
   IN2_i <= "00111001101000101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110111";
   IN2_i <= "01100111010010100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100111011";
   IN2_i <= "01111010001001100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110011110";
   IN2_i <= "00000100010001001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010110101";
   IN2_i <= "00101110011000010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001100100";
   IN2_i <= "00100101100010000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111011101";
   IN2_i <= "01110010011100111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000000010";
   IN2_i <= "00011011001011101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101110111";
   IN2_i <= "00111111111010010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111110000";
   IN2_i <= "00000010110011001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011100101";
   IN2_i <= "01111000000000100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011101";
   IN2_i <= "01101110011110011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010101";
   IN2_i <= "01011011001111110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110000111";
   IN2_i <= "00111101100111100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001100000";
   IN2_i <= "01010111011001000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001011";
   IN2_i <= "00011101100010101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010010000";
   IN2_i <= "01000110111111101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000101001";
   IN2_i <= "01110011111011101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010111000";
   IN2_i <= "00101101001000100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110001101";
   IN2_i <= "01000001110111000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000010011";
   IN2_i <= "00111111101010001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100011000";
   IN2_i <= "01010001101100110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100011100";
   IN2_i <= "01111111010010110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001010";
   IN2_i <= "01001000000001110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001010010";
   IN2_i <= "01001111010100111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010101011";
   IN2_i <= "01011101100010110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011101000";
   IN2_i <= "01111010000011111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001101000";
   IN2_i <= "00000011010010100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110001";
   IN2_i <= "01111100110000111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111001001";
   IN2_i <= "00001000011000100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010100110";
   IN2_i <= "01000011101110000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001001101";
   IN2_i <= "01111000111100110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010111010";
   IN2_i <= "01111101000110111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111000111";
   IN2_i <= "01110010111110101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010110110";
   IN2_i <= "01100101001100101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011001010";
   IN2_i <= "00001001100100101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001010110";
   IN2_i <= "01110101010011110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111010011";
   IN2_i <= "00101000110110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001101110";
   IN2_i <= "00110011011100101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001011001";
   IN2_i <= "01000001111010101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010010101";
   IN2_i <= "01001001010011111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010101001";
   IN2_i <= "01000001111011010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001101001";
   IN2_i <= "00111111011111001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011001100";
   IN2_i <= "00110111011110000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100110";
   IN2_i <= "00111010011111000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111001100";
   IN2_i <= "00001011100101011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011101110";
   IN2_i <= "01000011111100010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110001100";
   IN2_i <= "00111111111000010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101001001";
   IN2_i <= "00000010100001001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111010110";
   IN2_i <= "01101010111111111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010101000";
   IN2_i <= "01111010000001010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000011011";
   IN2_i <= "00001100101111011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110111101";
   IN2_i <= "00000111000010100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110000011";
   IN2_i <= "01001010010110000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011000";
   IN2_i <= "00011110011011110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111101010";
   IN2_i <= "01110101011010101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101110110";
   IN2_i <= "00000001011011110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100011010";
   IN2_i <= "00101110011100011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011110111";
   IN2_i <= "00100000100010111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111010001";
   IN2_i <= "00000100011110101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011101010";
   IN2_i <= "01110101000100101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001000110";
   IN2_i <= "01010110010101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100110111";
   IN2_i <= "01100010101001110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111000100";
   IN2_i <= "01011110000000110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010010101";
   IN2_i <= "01001101010001101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101010001";
   IN2_i <= "00110010000001010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101101110";
   IN2_i <= "01011101011001001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100100000";
   IN2_i <= "01000000100100101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000110101";
   IN2_i <= "01111111010111100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101011";
   IN2_i <= "00100101111011101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100110100";
   IN2_i <= "01100111011000011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100100100";
   IN2_i <= "01001100011010111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110100001";
   IN2_i <= "01001111111110011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001011001";
   IN2_i <= "00110111111100101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001010010";
   IN2_i <= "01010011111110100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001110011";
   IN2_i <= "00101010101100000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010010000";
   IN2_i <= "00101110011101000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110010101";
   IN2_i <= "00111111011110011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111011000";
   IN2_i <= "00000111010101010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010001100";
   IN2_i <= "01110111001001001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101111101";
   IN2_i <= "00100001011110110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001011111";
   IN2_i <= "00011110100001100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001101110";
   IN2_i <= "00101001100100110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011101011";
   IN2_i <= "00101000001010111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001110000";
   IN2_i <= "00000001111001011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011111000";
   IN2_i <= "00011111100110111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001001010";
   IN2_i <= "00110000100101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011001010";
   IN2_i <= "01101111011101110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110101110111";
   IN2_i <= "01001110000101001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101010011";
   IN2_i <= "00110110001001101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100100001";
   IN2_i <= "01111111000110110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110011101";
   IN2_i <= "00101010011111000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011010000";
   IN2_i <= "00111010100101011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100001001";
   IN2_i <= "00010100000001110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000101101";
   IN2_i <= "00100111001010101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111101";
   IN2_i <= "01111100111011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101011000";
   IN2_i <= "00011110011010001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001000110";
   IN2_i <= "01011100111000001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100001011";
   IN2_i <= "00001101001010000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010010100";
   IN2_i <= "01111110101100111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110010110";
   IN2_i <= "00000001011001111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001110010";
   IN2_i <= "01111100110011000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010010110";
   IN2_i <= "00100111111100101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100101111";
   IN2_i <= "00100110001010001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110001011";
   IN2_i <= "00110100000010011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101000";
   IN2_i <= "00011010111100100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110101101";
   IN2_i <= "00101101011101011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010011110";
   IN2_i <= "00010111010111100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010011111";
   IN2_i <= "00111110110101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101101111";
   IN2_i <= "01001010111110110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100000000";
   IN2_i <= "00100101000001000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100110101";
   IN2_i <= "00111011000100101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010000100";
   IN2_i <= "01000111011011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001110100";
   IN2_i <= "00001000010001100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100110110";
   IN2_i <= "01010101101010110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111000111";
   IN2_i <= "01001000010011111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001101101";
   IN2_i <= "01100001011110110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111010010";
   IN2_i <= "01000110001001111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011011000";
   IN2_i <= "01100100000111111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110001010";
   IN2_i <= "00111011011111010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000001011";
   IN2_i <= "00110101011011110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111111001111";
   IN2_i <= "00100101010101100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111011001";
   IN2_i <= "00010011001001110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101001";
   IN2_i <= "01000000111101101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010110111";
   IN2_i <= "01111000111111011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111110001";
   IN2_i <= "00011110011000011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011001";
   IN2_i <= "00010111101011110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100000111";
   IN2_i <= "01011010111000101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001101100";
   IN2_i <= "00011101110001000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101001110";
   IN2_i <= "01000100101101111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010101111";
   IN2_i <= "01111001111101101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101100110";
   IN2_i <= "00111111011110000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100110101";
   IN2_i <= "00100000100111001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010101100";
   IN2_i <= "01010111100100000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010011101";
   IN2_i <= "00110101111010001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001000101";
   IN2_i <= "01010011010110011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100001111";
   IN2_i <= "00000100011101000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000110101";
   IN2_i <= "01010011010111100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011011";
   IN2_i <= "00110111110001111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101111100";
   IN2_i <= "00001001100100010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000011111";
   IN2_i <= "01111010000111001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100100011";
   IN2_i <= "01000011010100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110001100";
   IN2_i <= "01011010100101011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100101011";
   IN2_i <= "01001011101001100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000101111";
   IN2_i <= "01101100000011001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101111101";
   IN2_i <= "01101100011110101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000011100";
   IN2_i <= "00111100000111100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111110100";
   IN2_i <= "01011001111010011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100001111";
   IN2_i <= "01010001011001110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101010";
   IN2_i <= "01011010100110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001100100";
   IN2_i <= "00100000000101100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010111111";
   IN2_i <= "01101010010110101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101100011";
   IN2_i <= "01111001011011101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111100101";
   IN2_i <= "01101010110001001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010101000";
   IN2_i <= "00001110000110101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010001010";
   IN2_i <= "01010111111101001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001011";
   IN2_i <= "01001110101011011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100100101";
   IN2_i <= "01011011110000111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011100111";
   IN2_i <= "00101101000100101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010010000";
   IN2_i <= "00001101000000101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101001110";
   IN2_i <= "00101111110001000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111010000";
   IN2_i <= "01010010000101000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111011011";
   IN2_i <= "00110000001011000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111011110";
   IN2_i <= "00110011010000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100011010";
   IN2_i <= "01111000011011001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010101110";
   IN2_i <= "01101101011011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101001100";
   IN2_i <= "00001100001011101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110001111";
   IN2_i <= "00010100010001000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100111100";
   IN2_i <= "00100001110100110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000001011";
   IN2_i <= "00010111011001001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101011";
   IN2_i <= "01000001110000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110111011";
   IN2_i <= "00011101011001111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011100000";
   IN2_i <= "00111001010101001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100100001";
   IN2_i <= "01001111100110110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100001110";
   IN2_i <= "00101011101001001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100111011";
   IN2_i <= "00111110001011011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111100100";
   IN2_i <= "01010110000010001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111111001";
   IN2_i <= "01111101011101110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111101010";
   IN2_i <= "00001110000011110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001011010";
   IN2_i <= "00011100000101101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011101011";
   IN2_i <= "00111111100000101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010101000";
   IN2_i <= "00010000000111101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110010111";
   IN2_i <= "00010110100100001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100010101";
   IN2_i <= "01000010001101100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010110011";
   IN2_i <= "01001011100110010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010100000";
   IN2_i <= "00110101111010101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111111001";
   IN2_i <= "01001000011101111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001000";
   IN2_i <= "01011010011111101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100110010";
   IN2_i <= "00111001001100010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101110100";
   IN2_i <= "01010111100111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001000110";
   IN2_i <= "01000111001110010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011000110";
   IN2_i <= "01111010011100101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011110110";
   IN2_i <= "01001101111100011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011111010";
   IN2_i <= "00010100110111110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001010010";
   IN2_i <= "01000110101011001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110101110";
   IN2_i <= "01100111001010110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001010100";
   IN2_i <= "00010100101101010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111100001";
   IN2_i <= "00111001100110111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001100001";
   IN2_i <= "01111101000110011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000110011";
   IN2_i <= "00000011101100011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011111010";
   IN2_i <= "00011000000001000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010111010";
   IN2_i <= "00011110110011011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111111101";
   IN2_i <= "01111100011000110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111111101";
   IN2_i <= "01100000000010000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000100110";
   IN2_i <= "01101000000111110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010000010";
   IN2_i <= "00011111010111101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111110";
   IN2_i <= "00001101000100000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101000010";
   IN2_i <= "00111011001100111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010010011";
   IN2_i <= "01100101010011101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000110010";
   IN2_i <= "00001101010011100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111011011";
   IN2_i <= "01011000001000110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101011001";
   IN2_i <= "01110010110001110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011011010";
   IN2_i <= "00001000110001011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101111011";
   IN2_i <= "00111001011010110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100010100";
   IN2_i <= "01100010101001000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010110100";
   IN2_i <= "01110101001111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010100110";
   IN2_i <= "00100010111000001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111101001";
   IN2_i <= "01101010101010101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100000001";
   IN2_i <= "01101000110100011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000100000";
   IN2_i <= "01010011000011110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001000101";
   IN2_i <= "01001000110011111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011011101";
   IN2_i <= "00111101000010110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111110001";
   IN2_i <= "01111011001001011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101101110";
   IN2_i <= "00011110111110111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101001110";
   IN2_i <= "01011010100101011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001011";
   IN2_i <= "00110000110011001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101011001";
   IN2_i <= "00001011000110101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011011011";
   IN2_i <= "01000011100011111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000111111";
   IN2_i <= "00110010101001010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111111111";
   IN2_i <= "01110010000000010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010011000";
   IN2_i <= "00101001000101001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010001110";
   IN2_i <= "00000100101110110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001100000";
   IN2_i <= "00100110110011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110101";
   IN2_i <= "00101001111111100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010010";
   IN2_i <= "01011111110100001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101001111";
   IN2_i <= "01101000011110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111100110";
   IN2_i <= "01110101011010001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000001110";
   IN2_i <= "01111111100000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010011000";
   IN2_i <= "00011000000100110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010011111";
   IN2_i <= "00001011110100001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001010000";
   IN2_i <= "00011001011110011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101110100";
   IN2_i <= "01001011001100010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100100011010";
   IN2_i <= "01011011100000100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101011001";
   IN2_i <= "01111110111010001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110000010";
   IN2_i <= "00011000101111111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001111000";
   IN2_i <= "01100110011100101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111011010";
   IN2_i <= "01101101100110110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010110";
   IN2_i <= "01011100100011100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101000111";
   IN2_i <= "01110010110100111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010011101";
   IN2_i <= "01101110110001010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001110010";
   IN2_i <= "01100010011000100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110110010";
   IN2_i <= "01011000101000111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110010010";
   IN2_i <= "00011011111101110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001010001";
   IN2_i <= "01110001110111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101001001";
   IN2_i <= "01111110001011001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000111110";
   IN2_i <= "00011011101110111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111011111";
   IN2_i <= "01001110010010010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000011100";
   IN2_i <= "01001110000101011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001000110";
   IN2_i <= "00100001101000011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101110";
   IN2_i <= "01010001010001100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100101001";
   IN2_i <= "01100001100100110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111010001";
   IN2_i <= "01100010110100000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100111110";
   IN2_i <= "01110110000000111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010011010";
   IN2_i <= "01111111111100100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010010001";
   IN2_i <= "01000010011000011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100101010";
   IN2_i <= "01100110110001111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001101010";
   IN2_i <= "00010000110000000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110101001";
   IN2_i <= "00111000101100111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100001110";
   IN2_i <= "00100000001010101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111000";
   IN2_i <= "00110000010100111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010110";
   IN2_i <= "00011000000001011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110000";
   IN2_i <= "00011010000001110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010110111";
   IN2_i <= "00010010101110111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010110100";
   IN2_i <= "00011011110000001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100001110";
   IN2_i <= "00001111010100110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110011100";
   IN2_i <= "00010011010001001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001011010";
   IN2_i <= "01110100011011100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110101101";
   IN2_i <= "00110111010011101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010111101";
   IN2_i <= "01100011000010011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111110100";
   IN2_i <= "01001010010001000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100100100";
   IN2_i <= "01011101111111111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011001011";
   IN2_i <= "00110010100001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111100000";
   IN2_i <= "01101101010101101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101110111";
   IN2_i <= "00010111110101101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000111101";
   IN2_i <= "01010111000111101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110101100";
   IN2_i <= "01111011000001110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110000111";
   IN2_i <= "00111110100001111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001010111";
   IN2_i <= "01001010000111110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001010010";
   IN2_i <= "00100100101110001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111010111";
   IN2_i <= "00110010001101000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001010100";
   IN2_i <= "00011011011100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100010100";
   IN2_i <= "01010110010100110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000000001";
   IN2_i <= "00110111010100111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101011000";
   IN2_i <= "01011000011000000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000010111";
   IN2_i <= "00100011010111101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100101011";
   IN2_i <= "01101001001000011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011001001";
   IN2_i <= "01111111001000101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011001000";
   IN2_i <= "00110111011100010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101000001";
   IN2_i <= "00100110111011101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110101010";
   IN2_i <= "01100000010010100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011011000";
   IN2_i <= "01000111011111101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000111010";
   IN2_i <= "00100101001011100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100010111";
   IN2_i <= "00111111100110011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010000100";
   IN2_i <= "00111011100101011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010101000";
   IN2_i <= "00000000000001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011100";
   IN2_i <= "01110011110111110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111010010";
   IN2_i <= "01101010111110100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000101110";
   IN2_i <= "00011110111000101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000110001";
   IN2_i <= "00010010100111100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100011001";
   IN2_i <= "00110101000111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100101111";
   IN2_i <= "00111111001000101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100111011";
   IN2_i <= "01111001010011010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101010110";
   IN2_i <= "01100101110010100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001010010";
   IN2_i <= "01001100011001101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110000000";
   IN2_i <= "01110101011111010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111111101";
   IN2_i <= "01011101011011110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001110000";
   IN2_i <= "01110001011011100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110010001";
   IN2_i <= "01001000000010100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000101100";
   IN2_i <= "01010011101110111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101101110";
   IN2_i <= "01011101000010111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010010101";
   IN2_i <= "01000101111001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101001011";
   IN2_i <= "01111011101111010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000001001";
   IN2_i <= "00001110001001100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101011101";
   IN2_i <= "01101111011111010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010001110";
   IN2_i <= "00100011110100010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101100011";
   IN2_i <= "01001111101001101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000100101";
   IN2_i <= "00000011110011101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101000010";
   IN2_i <= "01101000011011101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011001101";
   IN2_i <= "01011111100100000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011000011";
   IN2_i <= "00010100000001110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001100010";
   IN2_i <= "01110110100001010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101001100";
   IN2_i <= "01111010011101111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111111110";
   IN2_i <= "00010111001010000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110010111";
   IN2_i <= "01101101000011011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010111101";
   IN2_i <= "00011111101010111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010011101";
   IN2_i <= "00110010010010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110111";
   IN2_i <= "00101000110100001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100011111";
   IN2_i <= "00100111011011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101101010";
   IN2_i <= "00010000001000110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011000000";
   IN2_i <= "00100011011011100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001010101";
   IN2_i <= "00000101010001010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110011";
   IN2_i <= "00100101110000000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100100111";
   IN2_i <= "00010100101101010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011010011";
   IN2_i <= "00100011100110110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100010101";
   IN2_i <= "00001111010001100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001000010";
   IN2_i <= "00101001110100110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011110010";
   IN2_i <= "00100100101110111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000010000";
   IN2_i <= "00110001011011111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111101101";
   IN2_i <= "01001010100100010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011111101";
   IN2_i <= "00000111010000110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101001100";
   IN2_i <= "00001110101011110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111111010";
   IN2_i <= "01001001011001110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111011100";
   IN2_i <= "01010000101011000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101101110";
   IN2_i <= "01000110111101110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101001010";
   IN2_i <= "01100110001000111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010000111";
   IN2_i <= "00000011000010000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001001001";
   IN2_i <= "01010100011010101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100011001";
   IN2_i <= "01010110001000101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101111101";
   IN2_i <= "01010101000000110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110011010";
   IN2_i <= "01011110111110010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101001010";
   IN2_i <= "00001010100100010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100010110";
   IN2_i <= "00000111110110001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101000011";
   IN2_i <= "01101010100011001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010001011";
   IN2_i <= "00110100011010001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110001101";
   IN2_i <= "01000111000101010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001011011";
   IN2_i <= "00110101011100101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001101100";
   IN2_i <= "00000111001100111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100001100";
   IN2_i <= "01011010001001101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100101100";
   IN2_i <= "00111011100010000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111100011";
   IN2_i <= "00111110000111111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100100011";
   IN2_i <= "01100000011010000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011011010";
   IN2_i <= "00000011010010111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111111000";
   IN2_i <= "00010011001111111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000101110";
   IN2_i <= "00110111010011010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010011101";
   IN2_i <= "01100000010110101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111110101";
   IN2_i <= "00101000011001110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111010111";
   IN2_i <= "00001001000111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111101";
   IN2_i <= "00110100111111101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101011010";
   IN2_i <= "01100101110110000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011111111";
   IN2_i <= "00110011000011101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110110110";
   IN2_i <= "01000111110111010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100100111";
   IN2_i <= "01111110101100001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001111000";
   IN2_i <= "00010011001110100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110101101";
   IN2_i <= "01011011110011111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101111001";
   IN2_i <= "00101100101110100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100000011";
   IN2_i <= "01101101000000001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011000101";
   IN2_i <= "00111011100100011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111001010";
   IN2_i <= "00010010001011111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101000000";
   IN2_i <= "01001011011111110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010110110";
   IN2_i <= "00010000110110110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101110110";
   IN2_i <= "01100011011011111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010011";
   IN2_i <= "00111000011101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101111101";
   IN2_i <= "01111011000000110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101000000";
   IN2_i <= "00100000001101000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001101111";
   IN2_i <= "01000011101011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001110101";
   IN2_i <= "00011100010100000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111110101";
   IN2_i <= "01111101000001101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000100101";
   IN2_i <= "01111000010100001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100100011";
   IN2_i <= "00100011000111011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101010100";
   IN2_i <= "01010000111011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001010000";
   IN2_i <= "01111111111111000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111011000";
   IN2_i <= "00010111100111110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110001011";
   IN2_i <= "00010111100100001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010011111";
   IN2_i <= "00111100111110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110111011";
   IN2_i <= "00000111000000001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100111001";
   IN2_i <= "00001101100101010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011100011";
   IN2_i <= "00111110010000000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111111111";
   IN2_i <= "01111011101100001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000101011";
   IN2_i <= "01001011001101000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101010111";
   IN2_i <= "00010101110111011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111011100";
   IN2_i <= "01001101001100111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001001101";
   IN2_i <= "01101110110110101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010110000";
   IN2_i <= "01010011100101111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111111000";
   IN2_i <= "01000000111111100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110001111";
   IN2_i <= "01111110110000111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001010001";
   IN2_i <= "01101001011010100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010110010";
   IN2_i <= "00010101001111011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111010101";
   IN2_i <= "01101111000100100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101110001";
   IN2_i <= "01110001001010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000000000";
   IN2_i <= "01100101001110001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101000010";
   IN2_i <= "01010101110110000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001111010";
   IN2_i <= "01100011111100011";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110001111";
   IN2_i <= "00011110001000111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111000011";
   IN2_i <= "01100111001010001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110110010";
   IN2_i <= "00110011011101001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001010010";
   IN2_i <= "00100001001101010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011010110";
   IN2_i <= "01010000101011110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111011110";
   IN2_i <= "01010111101011010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001110111";
   IN2_i <= "00001011110110011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001100101";
   IN2_i <= "00011010110100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111010110";
   IN2_i <= "00000111110111010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001001000";
   IN2_i <= "01011000011111100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000010101";
   IN2_i <= "01100101000101100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011000010";
   IN2_i <= "00000110001011110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011100101";
   IN2_i <= "00101111110100100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111101010";
   IN2_i <= "01110000110111000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001101001";
   IN2_i <= "00001100010001001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111101000";
   IN2_i <= "01011011100010011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011111000";
   IN2_i <= "01011111001001001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111011010";
   IN2_i <= "00111111100001110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011001000";
   IN2_i <= "01011101101000101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011110101";
   IN2_i <= "01010101110111100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011111110";
   IN2_i <= "00000100001100010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000010110";
   IN2_i <= "01111000100000001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011110110";
   IN2_i <= "00101001011101100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101111";
   IN2_i <= "01100111011110010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100111010";
   IN2_i <= "01100111111101010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010110110";
   IN2_i <= "00000100011011110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001010";
   IN2_i <= "01111010011101111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101111111";
   IN2_i <= "01010111011100101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000101011";
   IN2_i <= "00110001010110010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100001011";
   IN2_i <= "01110000001110001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101000110";
   IN2_i <= "00101110110100111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010101011";
   IN2_i <= "01111001100111110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001101111";
   IN2_i <= "01000011011010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001111110";
   IN2_i <= "00100000011110000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011100001";
   IN2_i <= "00100000010011010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000000001";
   IN2_i <= "00000001111001001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001011100";
   IN2_i <= "00101100111101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011101100";
   IN2_i <= "00011101001111100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100011010";
   IN2_i <= "00100001001101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001110";
   IN2_i <= "00101000101101001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100100110";
   IN2_i <= "00101001010100000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011110010";
   IN2_i <= "00111110101011111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010001110";
   IN2_i <= "00010011000011111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001110000";
   IN2_i <= "00010011001100101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000011000";
   IN2_i <= "00110101010000101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111001000";
   IN2_i <= "01111100100011010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111100101";
   IN2_i <= "01010000001010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010110010";
   IN2_i <= "01110110110001000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111000111";
   IN2_i <= "01101000100101100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001001111";
   IN2_i <= "01011000101101110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110100011";
   IN2_i <= "00111101101000110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110111011";
   IN2_i <= "01110011110101000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001111100";
   IN2_i <= "01011110011100011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010011010";
   IN2_i <= "00100000111101101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111111000";
   IN2_i <= "01111110111101101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001000000";
   IN2_i <= "01000110000111110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000101111";
   IN2_i <= "00011011001101010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010111000";
   IN2_i <= "00001101011110100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101100111";
   IN2_i <= "01110011101000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100111000";
   IN2_i <= "01101110101111111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110100100";
   IN2_i <= "01100101100011000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101000010";
   IN2_i <= "00100010101101000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100001110";
   IN2_i <= "01100000101110110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010101110";
   IN2_i <= "00010000000111110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001110001";
   IN2_i <= "01101111001111110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100101000";
   IN2_i <= "01001011000000001";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011110110";
   IN2_i <= "01000011010111010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100010101";
   IN2_i <= "01101011100010110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011000110111";
   IN2_i <= "01000111010110010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111001011";
   IN2_i <= "00111011101011110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001011101";
   IN2_i <= "00100111011101010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001101100";
   IN2_i <= "00110010100011110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010001100";
   IN2_i <= "01011111111100110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000100101";
   IN2_i <= "01110011001111010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101011010";
   IN2_i <= "00011011010111110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100100011";
   IN2_i <= "00100000111011000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011010010";
   IN2_i <= "01101100000010100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110101010";
   IN2_i <= "00001110001010110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111111111";
   IN2_i <= "00011101011110110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100011100";
   IN2_i <= "01111000001001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001101001";
   IN2_i <= "01111001101011000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111011100";
   IN2_i <= "01011100011111000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111101011";
   IN2_i <= "00010010110101001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111011110";
   IN2_i <= "01110101110001011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110010010";
   IN2_i <= "01001110001011110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000100001";
   IN2_i <= "00001100101100011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010110011";
   IN2_i <= "01111101000000010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100111";
   IN2_i <= "00100100111010010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010101000110";
   IN2_i <= "00010010001111100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111010110";
   IN2_i <= "01110000000000100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110111110101";
   IN2_i <= "00110001010111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110101011";
   IN2_i <= "00010111010001100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001100100";
   IN2_i <= "01110000001001101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010010100";
   IN2_i <= "00011010011010000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100001000";
   IN2_i <= "00100001111010110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011010110";
   IN2_i <= "00100111110101001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101001101";
   IN2_i <= "01111100010101111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100000010";
   IN2_i <= "00000011110100010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101010";
   IN2_i <= "00111000010101110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111001";
   IN2_i <= "01110011010000001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111100";
   IN2_i <= "00100110100100010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100100100";
   IN2_i <= "00011001000001001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100010101";
   IN2_i <= "01010101101011101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110001011";
   IN2_i <= "00110011111111010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110011";
   IN2_i <= "01011110011110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000101110";
   IN2_i <= "00000001110000011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000100101";
   IN2_i <= "01110100110011001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100011001";
   IN2_i <= "00111000000110110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101110101";
   IN2_i <= "00010110110100000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110011111";
   IN2_i <= "00110111100000000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010011100";
   IN2_i <= "00011000000100001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100101";
   IN2_i <= "01101001010001110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000110010";
   IN2_i <= "00100110011011101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011100010";
   IN2_i <= "00011111001111011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001001101";
   IN2_i <= "01001011000001100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101111011";
   IN2_i <= "00100010011010110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110110";
   IN2_i <= "00100001011010001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111000011";
   IN2_i <= "01100011011111001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101010000";
   IN2_i <= "01111101111010110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111011110";
   IN2_i <= "01110000011101111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001101010";
   IN2_i <= "00110010011000011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111001101";
   IN2_i <= "00001111111011000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100010111";
   IN2_i <= "01010001000100100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000001010";
   IN2_i <= "01111110100110101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111110000";
   IN2_i <= "01011111011010001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011000010";
   IN2_i <= "01001101001100111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001110010";
   IN2_i <= "00111101001011110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000000101";
   IN2_i <= "00101000010011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101101101";
   IN2_i <= "00110111101011111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001011110";
   IN2_i <= "01000000011010000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001010001";
   IN2_i <= "00101101010010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011001";
   IN2_i <= "01010101101001010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110000011";
   IN2_i <= "01000110101100001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011101100";
   IN2_i <= "01100011101101010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100100000";
   IN2_i <= "00101011010001011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111001010";
   IN2_i <= "01001101101110101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000011101";
   IN2_i <= "00110100101101001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001101111";
   IN2_i <= "01101100011111101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100000100";
   IN2_i <= "00001100110100100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110101100";
   IN2_i <= "01010001111000111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001000010";
   IN2_i <= "01110010101010110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000000101";
   IN2_i <= "00100100011000001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010010";
   IN2_i <= "00011001110001111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011011";
   IN2_i <= "01110100110110010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011111000";
   IN2_i <= "01000100000010100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010111100";
   IN2_i <= "01111111101111000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000010000";
   IN2_i <= "01100001101010100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011011101";
   IN2_i <= "00011001001000101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111100100";
   IN2_i <= "01001010110100110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100110000";
   IN2_i <= "01111111000100001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001010101";
   IN2_i <= "00001001100110010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011110100";
   IN2_i <= "00101000111100010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010100";
   IN2_i <= "00101110100100100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101110001";
   IN2_i <= "01111011110001001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110100111";
   IN2_i <= "00000100011111110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011110000";
   IN2_i <= "01011100111100100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010100111";
   IN2_i <= "00101001000100100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101010111";
   IN2_i <= "00000010100011110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111111000";
   IN2_i <= "01101110111010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011100110";
   IN2_i <= "01100011111110001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011110101";
   IN2_i <= "01001010000111011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110000000";
   IN2_i <= "00010111110001111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101100010";
   IN2_i <= "00010101111010011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011110010";
   IN2_i <= "00011111010011001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000111100";
   IN2_i <= "00000001001101010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010100111";
   IN2_i <= "00010011100001001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100000000";
   IN2_i <= "00100001100001000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100001111";
   IN2_i <= "01101110000101011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011001010";
   IN2_i <= "01111110110000001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011011000";
   IN2_i <= "00111011101101000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101100000";
   IN2_i <= "00111010000100011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010011010";
   IN2_i <= "01010000101010100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001011110";
   IN2_i <= "01001111100001100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001010101";
   IN2_i <= "01100010010010011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010100010";
   IN2_i <= "00111101100000010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101001";
   IN2_i <= "01011011001111011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110100010";
   IN2_i <= "01111100110010101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101010011";
   IN2_i <= "00110101010111101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010000";
   IN2_i <= "01001101011101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001101101";
   IN2_i <= "01111000011101010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001001010";
   IN2_i <= "01100011000111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001011111";
   IN2_i <= "01000110110110111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011010101";
   IN2_i <= "00001011100110011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111001011";
   IN2_i <= "01101010001011100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100100000";
   IN2_i <= "00010100000111111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110001101";
   IN2_i <= "01110010101101100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011111";
   IN2_i <= "00101100000001000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111000001";
   IN2_i <= "01101010000001010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101100101";
   IN2_i <= "01010001010111111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010110011";
   IN2_i <= "00000110100110101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000101001";
   IN2_i <= "01011011100100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001110100";
   IN2_i <= "01111000100110000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010000001";
   IN2_i <= "00111000000101111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100101010";
   IN2_i <= "00010101101000011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110101011";
   IN2_i <= "00010100110011110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100110010";
   IN2_i <= "01001111100011111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110110000";
   IN2_i <= "01000010010011111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111011110";
   IN2_i <= "01011111011111000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101111011";
   IN2_i <= "01001111110111000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111101000";
   IN2_i <= "01111101011011101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101111110";
   IN2_i <= "00101101001000001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111110000";
   IN2_i <= "01111100000000111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000110110";
   IN2_i <= "01111110111101000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001000000";
   IN2_i <= "01101000101011010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000011011";
   IN2_i <= "00000100010111100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000101100";
   IN2_i <= "00010110001110001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000001100";
   IN2_i <= "00001100111010111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100101110";
   IN2_i <= "00001001101110001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101001000";
   IN2_i <= "00111011110111010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110011110";
   IN2_i <= "00100110010101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101011";
   IN2_i <= "01001010111000110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101101001";
   IN2_i <= "01000111001011101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001101";
   IN2_i <= "00111101111010111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110010011";
   IN2_i <= "00000110001010001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000011111";
   IN2_i <= "01101010011110001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010101011";
   IN2_i <= "01000010100101011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100100110";
   IN2_i <= "00101011111100010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111000100";
   IN2_i <= "01101010101110010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000100011";
   IN2_i <= "00010010101110011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011010001";
   IN2_i <= "01011100101101010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110110001";
   IN2_i <= "01010100000111101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000101";
   IN2_i <= "01000000111011101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001000011";
   IN2_i <= "01001001100010110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111100001";
   IN2_i <= "00111110001011010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100101111";
   IN2_i <= "00110101010001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111101110";
   IN2_i <= "01111011001010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001101000";
   IN2_i <= "01011011000010111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101001001";
   IN2_i <= "01010001010011101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001001011";
   IN2_i <= "01100101011110011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101101000";
   IN2_i <= "01100000000101110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001101001";
   IN2_i <= "00001000111111010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110111100";
   IN2_i <= "01001100100000110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101001101";
   IN2_i <= "00010001100010010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000100101";
   IN2_i <= "00011111110000001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000000110";
   IN2_i <= "01010111011111011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101101111";
   IN2_i <= "01000010011110000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110011110";
   IN2_i <= "01011001000010001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110101011";
   IN2_i <= "01101110101001000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010111001";
   IN2_i <= "00011101110110010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000110";
   IN2_i <= "01111000100111111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111000111";
   IN2_i <= "00011001010110001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100010000";
   IN2_i <= "01111100001111110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011101001";
   IN2_i <= "01000011100111110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001000000";
   IN2_i <= "00111111101010101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100000100";
   IN2_i <= "01000101100111000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000101000";
   IN2_i <= "00111100000001101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000000001";
   IN2_i <= "00111111011010101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010110";
   IN2_i <= "00111001111100101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010111011";
   IN2_i <= "00011111101011110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011101001";
   IN2_i <= "01110001111010000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101101111";
   IN2_i <= "01011000110101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001011010";
   IN2_i <= "01110100110100101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101011";
   IN2_i <= "00010101000101011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010100100";
   IN2_i <= "01101001110011000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011111101";
   IN2_i <= "01000000111000000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100010000";
   IN2_i <= "00001011010001000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010110010";
   IN2_i <= "00101100010110001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111101000";
   IN2_i <= "00101000101101111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100100001";
   IN2_i <= "01011011011101010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000101110";
   IN2_i <= "01110001110011011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010000011";
   IN2_i <= "00011111101101110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110110000";
   IN2_i <= "00110100101001000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101001100";
   IN2_i <= "00101001011010011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111011111";
   IN2_i <= "01101101111001100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100110111";
   IN2_i <= "01001001000111100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001111001";
   IN2_i <= "00001001001101101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100101111";
   IN2_i <= "00001000010100110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100011001";
   IN2_i <= "00100000011101001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011110";
   IN2_i <= "00000111111111001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011010101";
   IN2_i <= "01010100111111011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100111001";
   IN2_i <= "00010000011110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000110100";
   IN2_i <= "01101001111001100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001111";
   IN2_i <= "00010001011011010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000111101";
   IN2_i <= "00010111100101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010011000";
   IN2_i <= "00000010110110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110110010";
   IN2_i <= "01111111000101111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011111101";
   IN2_i <= "00000100000011000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001100011";
   IN2_i <= "00110101101101111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001001101";
   IN2_i <= "00100010000110100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101111111";
   IN2_i <= "01111100100011011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100001001";
   IN2_i <= "01011010001110100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110100010";
   IN2_i <= "00000010001000011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010000100";
   IN2_i <= "01010100110010001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001111001";
   IN2_i <= "00010011011101100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000101010";
   IN2_i <= "01000101111100110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110111110";
   IN2_i <= "01111100010000010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111111111";
   IN2_i <= "01110010011010110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011111011";
   IN2_i <= "01110000011001111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111101110";
   IN2_i <= "01100011100101110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000110010";
   IN2_i <= "00111000100001001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101101001";
   IN2_i <= "00001110100110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000111101";
   IN2_i <= "00001100101111101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010111010";
   IN2_i <= "01010011011001100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100110100";
   IN2_i <= "00101110101011000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111110111";
   IN2_i <= "00000111010111000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110100100";
   IN2_i <= "00000100111000101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000010110";
   IN2_i <= "01111111000100010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100100100";
   IN2_i <= "00101110101001101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110100001";
   IN2_i <= "01110000110010100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100000111";
   IN2_i <= "01000001111100100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101111010";
   IN2_i <= "01000010000101001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000011000";
   IN2_i <= "00010101110001111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010110001";
   IN2_i <= "00110110011011011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110101";
   IN2_i <= "01100011011010000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011101001";
   IN2_i <= "01111001011101011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000100100";
   IN2_i <= "01001010100010110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001010010";
   IN2_i <= "00001000011101111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011011111";
   IN2_i <= "00100010010011011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010101";
   IN2_i <= "01110100100101000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110010110";
   IN2_i <= "00000111101101110";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100010110";
   IN2_i <= "01100101010110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100100101";
   IN2_i <= "00110000000001000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010111000";
   IN2_i <= "01010000111011110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101000";
   IN2_i <= "01100011001101101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101010010";
   IN2_i <= "00000101111010100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100101110";
   IN2_i <= "00010101111110101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100000011";
   IN2_i <= "01100111010001100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110011100";
   IN2_i <= "01010101001010111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001001010";
   IN2_i <= "00001111010011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101110101";
   IN2_i <= "01110011000011010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101101001";
   IN2_i <= "01110001011100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111111";
   IN2_i <= "00100011010011001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100100000";
   IN2_i <= "01110100011010100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101101010";
   IN2_i <= "00001110100110011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001001010";
   IN2_i <= "00110101101000101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110001100";
   IN2_i <= "00000011001101101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000011111";
   IN2_i <= "00010100000100100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100111101";
   IN2_i <= "00010011001100011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001111010";
   IN2_i <= "00010111000111001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111000001";
   IN2_i <= "01111000101100011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001001100001";
   IN2_i <= "00010000010001111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101010101";
   IN2_i <= "01001101111110110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010000100";
   IN2_i <= "00111000011101101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000000111";
   IN2_i <= "01000001111110001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010111000";
   IN2_i <= "00111110011011010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011000000";
   IN2_i <= "01000101011010010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011100101";
   IN2_i <= "00111011100001000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001001001";
   IN2_i <= "00001011110100110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111001001";
   IN2_i <= "01010010010010101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011110011";
   IN2_i <= "00111000110110101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110101110";
   IN2_i <= "00010110011100111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011100111";
   IN2_i <= "01011111100011000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110001010";
   IN2_i <= "00111011000011010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100100010";
   IN2_i <= "01000110010100011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111110000";
   IN2_i <= "00001110011100111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001111101";
   IN2_i <= "01010001101000001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101000111";
   IN2_i <= "00100000110100011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101100111";
   IN2_i <= "00100011010001010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100111000";
   IN2_i <= "00001000000101110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010111111";
   IN2_i <= "01101111101001101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000100111";
   IN2_i <= "00001011010101010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000011";
   IN2_i <= "01000010110111001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000110101";
   IN2_i <= "00110001010100000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100100111";
   IN2_i <= "01100111101001111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110010011";
   IN2_i <= "00101000000111010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110110000";
   IN2_i <= "01100001111011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010000010";
   IN2_i <= "01011111010010101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000111110";
   IN2_i <= "01100011001011111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101111110";
   IN2_i <= "01010111111111001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110101";
   IN2_i <= "00101110100100111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101110010";
   IN2_i <= "00101011011000110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001101110";
   IN2_i <= "00010101001011111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011000101";
   IN2_i <= "01000100100011001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111000110";
   IN2_i <= "01010010001101000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001011";
   IN2_i <= "01101101001110111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001101100";
   IN2_i <= "00110001001110011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001000110";
   IN2_i <= "00011111011110101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100110000";
   IN2_i <= "01100011010010110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010000100111";
   IN2_i <= "01111001010001110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000001101";
   IN2_i <= "01110011111010001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100000";
   IN2_i <= "01011100111100101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010001110";
   IN2_i <= "01000101111001011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001001";
   IN2_i <= "00011001101101011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100010111";
   IN2_i <= "01110101100010100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011101101";
   IN2_i <= "00001110010001110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101000";
   IN2_i <= "01010111110010110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101110111";
   IN2_i <= "00111100010001001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001101001";
   IN2_i <= "01100101101100110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001101010";
   IN2_i <= "01001011011011000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111100100";
   IN2_i <= "01101000010000011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000000";
   IN2_i <= "00001011010111000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100111101";
   IN2_i <= "01101010011011010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001100010";
   IN2_i <= "01011100101011000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011001011";
   IN2_i <= "00001001011111101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110110011";
   IN2_i <= "00000111010111011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001110100000";
   IN2_i <= "01011101110010101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101000100";
   IN2_i <= "00010001110000010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001100010";
   IN2_i <= "01001000011001100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101101100";
   IN2_i <= "00111010001000010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111000010";
   IN2_i <= "01011010101000110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010000101";
   IN2_i <= "01010010010100011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110001111";
   IN2_i <= "00011111001000000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010100000";
   IN2_i <= "00100101111101001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000111010";
   IN2_i <= "01111101000011001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100000010";
   IN2_i <= "01001011110110011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001101000";
   IN2_i <= "01111111101011101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101000110";
   IN2_i <= "01001110111101101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111010111";
   IN2_i <= "01001010011000000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011111110";
   IN2_i <= "01101011001001110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101000011";
   IN2_i <= "00101010011110110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100101";
   IN2_i <= "00000001011000010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011001";
   IN2_i <= "01011011001011011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000001001";
   IN2_i <= "00101110111100100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000100110";
   IN2_i <= "00010101101101001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010001101";
   IN2_i <= "01000111110100010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010011111";
   IN2_i <= "00111001101001111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101011000";
   IN2_i <= "00100011010010001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011000101";
   IN2_i <= "01111001111011110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000111000";
   IN2_i <= "01001100000010010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010001011";
   IN2_i <= "01101000100101000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011100111";
   IN2_i <= "01100001100010000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000100011";
   IN2_i <= "01010110000000111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110110111";
   IN2_i <= "00010000101010100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000000111";
   IN2_i <= "01000101101011010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010111010";
   IN2_i <= "01000000000110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100111101";
   IN2_i <= "00011011111010110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001011110";
   IN2_i <= "01110101100011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011111011";
   IN2_i <= "01111110010000011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100000010";
   IN2_i <= "00001011001000100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101001001";
   IN2_i <= "01000000000011111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110110010";
   IN2_i <= "00101101111110011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001011110";
   IN2_i <= "00000100111110101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110001110";
   IN2_i <= "01101011000111110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101001101";
   IN2_i <= "01011000010000101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111011110";
   IN2_i <= "00000010000100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111111001";
   IN2_i <= "00101011010101101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010101001";
   IN2_i <= "01010010010011101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110001000";
   IN2_i <= "01100010100011011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111011111";
   IN2_i <= "00000011010000001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111110111";
   IN2_i <= "01101011100011001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111101100";
   IN2_i <= "00110110111100001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010110100";
   IN2_i <= "00000001000001111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110000010";
   IN2_i <= "00011011111101110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000110000";
   IN2_i <= "00000001010010010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001111100";
   IN2_i <= "01000010010011101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011100011";
   IN2_i <= "01110111000000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011111100";
   IN2_i <= "01100011110000010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100100111";
   IN2_i <= "00001000110001101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010101111";
   IN2_i <= "00100001010010110";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000001000";
   IN2_i <= "00100110011001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000011001111";
   IN2_i <= "01001101010101110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110010010";
   IN2_i <= "01101101101010000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011100011";
   IN2_i <= "00010000110000111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110111000";
   IN2_i <= "01001110001100110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100001";
   IN2_i <= "01010000011110000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001111011";
   IN2_i <= "00101100101000001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000110100";
   IN2_i <= "00100001011111100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111100011";
   IN2_i <= "01101101100011100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110100010110";
   IN2_i <= "01000000111101101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010111010";
   IN2_i <= "01010110110011000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010101000";
   IN2_i <= "00110100110111000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110111010";
   IN2_i <= "01010011011100101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100001101";
   IN2_i <= "01000111000001011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000100001111";
   IN2_i <= "01011001000111011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110001111";
   IN2_i <= "00000011101011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011010011";
   IN2_i <= "01110101001111011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100111000";
   IN2_i <= "00000100001110100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100000011";
   IN2_i <= "00000111001001110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101100100";
   IN2_i <= "01001010000010111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101000000";
   IN2_i <= "00000010001000100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110011000";
   IN2_i <= "01111111010100110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111100000";
   IN2_i <= "01111000010110111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100001100";
   IN2_i <= "00001010100011000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100001111";
   IN2_i <= "00011000100010100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000101110";
   IN2_i <= "00100010111011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100010111";
   IN2_i <= "01100110100110100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001111001";
   IN2_i <= "00101000000110110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011001100";
   IN2_i <= "01111100110100101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001010100";
   IN2_i <= "01001011011011110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100011001";
   IN2_i <= "00111001100010000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000101110";
   IN2_i <= "00001010000101010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001100100";
   IN2_i <= "00000110101101011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001100110";
   IN2_i <= "00011000010000101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111100100";
   IN2_i <= "01000111100100100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011110100";
   IN2_i <= "00111000100010101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010100100";
   IN2_i <= "01110001111000101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100011011";
   IN2_i <= "00010110100001100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010101100";
   IN2_i <= "00011011101111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101101010";
   IN2_i <= "01111010001110010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101110110";
   IN2_i <= "01101101110100111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100101001";
   IN2_i <= "00111110100111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111010010";
   IN2_i <= "01101111100100011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101100011";
   IN2_i <= "00110100100101110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111001101";
   IN2_i <= "01101101111110111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111000";
   IN2_i <= "01000000011011110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010100";
   IN2_i <= "00110110111011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101111001";
   IN2_i <= "01011001010001100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110000010";
   IN2_i <= "00101100111110001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001101001";
   IN2_i <= "00010101111110100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010101111";
   IN2_i <= "01111010001001111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111111001";
   IN2_i <= "00111011010011011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000111100";
   IN2_i <= "01010111000010101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010011000";
   IN2_i <= "00001101101111000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001111011";
   IN2_i <= "00000101000111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001001010";
   IN2_i <= "00101010110000101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001110100";
   IN2_i <= "01101001010100000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111111011";
   IN2_i <= "01001010011100101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100010100";
   IN2_i <= "00011100111101010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100011101";
   IN2_i <= "00110100100000011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100111110";
   IN2_i <= "01000000010100101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011001101";
   IN2_i <= "01000100111100010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111011110";
   IN2_i <= "01000100000100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110010";
   IN2_i <= "00101001011010101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110010010";
   IN2_i <= "00110000010110111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110010100";
   IN2_i <= "01100011111100111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001111110";
   IN2_i <= "01100001011111101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111100010";
   IN2_i <= "00011011101101100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110101111";
   IN2_i <= "01010110011100111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011011111";
   IN2_i <= "01111110010110010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000010111";
   IN2_i <= "01100000010111011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011010001";
   IN2_i <= "00100010110011011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000110001";
   IN2_i <= "01101100110000011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000011011";
   IN2_i <= "01000000010110001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111010000";
   IN2_i <= "01000110111100111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001101110";
   IN2_i <= "00101001000101010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000100001";
   IN2_i <= "00111101110111001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110001000";
   IN2_i <= "01100000011110110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010101000";
   IN2_i <= "01000010100111011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101011100";
   IN2_i <= "01100111111100100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001110001";
   IN2_i <= "00100001101111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111111";
   IN2_i <= "01111001010010011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000010111";
   IN2_i <= "01100111101101111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110010101";
   IN2_i <= "00000011001100011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110011010";
   IN2_i <= "00010000110100001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110000010";
   IN2_i <= "00001100100001010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111011101";
   IN2_i <= "01011001000110011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000101101";
   IN2_i <= "00001000110110111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101101000";
   IN2_i <= "01011110011111001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100011";
   IN2_i <= "00010100000101111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000100010";
   IN2_i <= "01010001001110011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100011";
   IN2_i <= "00001010101010001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001010101";
   IN2_i <= "00101001101001010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110001";
   IN2_i <= "00010100101101000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110100110";
   IN2_i <= "01111111111100100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111001001";
   IN2_i <= "00011011100101110";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100111000";
   IN2_i <= "00100001001111000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010011010";
   IN2_i <= "01100000110001110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001101100";
   IN2_i <= "00110000011001101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011110101";
   IN2_i <= "00000001110011110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100001111";
   IN2_i <= "00100111010110010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010010110";
   IN2_i <= "01110001010110110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001010111";
   IN2_i <= "01011011001100001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011110100";
   IN2_i <= "00000001101000011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110011010";
   IN2_i <= "00010001101100110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100000100";
   IN2_i <= "01111011010010101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100011111";
   IN2_i <= "01010010010111010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000010111";
   IN2_i <= "00110001001011011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001111011";
   IN2_i <= "01010111111011001";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110001000";
   IN2_i <= "00101010111011001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000011111";
   IN2_i <= "01100010011001011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100100110";
   IN2_i <= "01001010001011100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001110111";
   IN2_i <= "01101010110101001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011011100";
   IN2_i <= "01011100000101000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011100001";
   IN2_i <= "01001101001001001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100100011";
   IN2_i <= "01110100111001111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001011110";
   IN2_i <= "01010001000001001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100010001";
   IN2_i <= "01010011101111011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010111";
   IN2_i <= "01001000001110101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010111111";
   IN2_i <= "00100111010111011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000101011";
   IN2_i <= "01100011110111011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000111000";
   IN2_i <= "00100011111111100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000111101";
   IN2_i <= "00101111101101010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111000101";
   IN2_i <= "01011110111101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000001110";
   IN2_i <= "00110000101101101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110000110";
   IN2_i <= "01101011100001011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101101001";
   IN2_i <= "01100111010011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000001010";
   IN2_i <= "00100010001101001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010101101";
   IN2_i <= "00111010101101010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111010001";
   IN2_i <= "01001110101001110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100011001";
   IN2_i <= "00111110110100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001101000";
   IN2_i <= "00010000110001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101011101";
   IN2_i <= "00111001101011101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000101111";
   IN2_i <= "01000011000001000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011100101";
   IN2_i <= "01010000111010100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110101001";
   IN2_i <= "01101111010110110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001110110";
   IN2_i <= "01011111110101111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110001110";
   IN2_i <= "00100000011111110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101101000";
   IN2_i <= "00100100100010101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111000110";
   IN2_i <= "01110101010000011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011101110";
   IN2_i <= "01110100000101100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110101111";
   IN2_i <= "01100100001011101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100011000";
   IN2_i <= "00100011001101111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101000000";
   IN2_i <= "00101010000011111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001000100";
   IN2_i <= "00001001101001001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011110010";
   IN2_i <= "00011111000010101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101011000";
   IN2_i <= "00011011101100111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010111011";
   IN2_i <= "01100001101110111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101100110";
   IN2_i <= "00100111000001111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000001011001";
   IN2_i <= "00000110001011010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111011010";
   IN2_i <= "01001110001011100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111100101";
   IN2_i <= "00000111000000111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110011111";
   IN2_i <= "01111011100000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110000000";
   IN2_i <= "01000110101010001";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100011010";
   IN2_i <= "01001100010110000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011111010";
   IN2_i <= "00000000011111010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100011101";
   IN2_i <= "00001100110001011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110000001";
   IN2_i <= "00111000001000000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011000110";
   IN2_i <= "01101110110011010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101111110";
   IN2_i <= "01111101110001100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101100010";
   IN2_i <= "00000001010111111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011000000";
   IN2_i <= "00000010100111011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100000";
   IN2_i <= "01111101110000001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100101011";
   IN2_i <= "01111111000010110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001111100";
   IN2_i <= "00100100101011111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101001100";
   IN2_i <= "00100100110001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010010110";
   IN2_i <= "01100111011110100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010100";
   IN2_i <= "00100110110011010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011000100";
   IN2_i <= "00110010001001110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111101";
   IN2_i <= "01000101111011011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011001010";
   IN2_i <= "01111101110110110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011100101";
   IN2_i <= "00000001010000010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110000111";
   IN2_i <= "00101001100101000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010101100";
   IN2_i <= "00011011111100110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011001110";
   IN2_i <= "00111011110101001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111100";
   IN2_i <= "00101111100100000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001001111";
   IN2_i <= "01011110000100111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111010010";
   IN2_i <= "00110011100000010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000000001";
   IN2_i <= "01010011001011110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000001000";
   IN2_i <= "00001011101101010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110111000";
   IN2_i <= "01010010100001001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011000101010";
   IN2_i <= "01101101101011001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100011011";
   IN2_i <= "01001010011010010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001001100";
   IN2_i <= "01001101110111100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110110001";
   IN2_i <= "00111010100100001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110110011";
   IN2_i <= "01001101010110001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000001100";
   IN2_i <= "01111010111101100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111111110";
   IN2_i <= "01001101110111011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101010110";
   IN2_i <= "00110101011010111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110100000";
   IN2_i <= "00001110010000010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000011101";
   IN2_i <= "00111111100011011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111001010";
   IN2_i <= "01111101110011100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111010100";
   IN2_i <= "00101101010010111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010001101010";
   IN2_i <= "00011110100100010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011101111000";
   IN2_i <= "01110100000000001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110111011";
   IN2_i <= "01011111111100111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100000110";
   IN2_i <= "01111011001011111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100001101";
   IN2_i <= "01111111001011111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010001010";
   IN2_i <= "00111000100011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101111101";
   IN2_i <= "01110001000110011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010001";
   IN2_i <= "00101101110100010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001000011";
   IN2_i <= "00011001011110100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110010100";
   IN2_i <= "01000010110001100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111010111";
   IN2_i <= "01011110110000000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011111001";
   IN2_i <= "01100010001111110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101110000";
   IN2_i <= "01101111111100111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000010100";
   IN2_i <= "00010001100100000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100110111110";
   IN2_i <= "01000100110110011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011101101";
   IN2_i <= "00101110101010110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011011101";
   IN2_i <= "00010100111011011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100000000";
   IN2_i <= "01100101001001000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110001001";
   IN2_i <= "01000111111111110";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101101101";
   IN2_i <= "00001110001001010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111110010";
   IN2_i <= "00001001110001010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101001111";
   IN2_i <= "00101001000001011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110011110";
   IN2_i <= "00111110011011110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101100110";
   IN2_i <= "00100100011101001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110010011";
   IN2_i <= "00111011110001111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010111010";
   IN2_i <= "00101000110010010";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000110110";
   IN2_i <= "01110000110010001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011100";
   IN2_i <= "00111100101011000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110111001";
   IN2_i <= "00011000101000111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110000011";
   IN2_i <= "01101001111110011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011100";
   IN2_i <= "01100011010100100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011100110";
   IN2_i <= "01001000100001111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100101010";
   IN2_i <= "00111110000010011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011110111";
   IN2_i <= "00010110100011111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100110000";
   IN2_i <= "00101000001010100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001110101";
   IN2_i <= "01000110111000010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111001001";
   IN2_i <= "00101101001011111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111111100";
   IN2_i <= "01100011101011010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010001101";
   IN2_i <= "01110100111000001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100110000";
   IN2_i <= "00111101110000111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101100110";
   IN2_i <= "01110100110111110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000000100";
   IN2_i <= "00010001100101110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110001";
   IN2_i <= "01001001011001101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100001001";
   IN2_i <= "01100011110001111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110011100";
   IN2_i <= "01000011000111000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010101111";
   IN2_i <= "01000100111010111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101011111";
   IN2_i <= "00111101010011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001011";
   IN2_i <= "00101100110111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001100001";
   IN2_i <= "01100001011001001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100011001";
   IN2_i <= "01000001000111110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100001011";
   IN2_i <= "01011100101110111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011011001";
   IN2_i <= "00011000111100000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000110000";
   IN2_i <= "00110111101011111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101111100";
   IN2_i <= "00001110101000000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001010111";
   IN2_i <= "01110001100100000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001110";
   IN2_i <= "00110111001001010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010011";
   IN2_i <= "00010000111010111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010111011101";
   IN2_i <= "01100110010101111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000011110";
   IN2_i <= "00000010011000100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100001000";
   IN2_i <= "01001010000010011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100110010";
   IN2_i <= "01110010001101110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000111011";
   IN2_i <= "01111010100110000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010011111";
   IN2_i <= "00111010111111110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001100110";
   IN2_i <= "00011010110111010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010001";
   IN2_i <= "01100010010001101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110010100";
   IN2_i <= "00010100000101010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010010110";
   IN2_i <= "01010010100001001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111110001";
   IN2_i <= "01100001000111110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111100111011";
   IN2_i <= "00010111011100101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001000010";
   IN2_i <= "01011010011010011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110101101";
   IN2_i <= "00101100010110011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101111100";
   IN2_i <= "01011100001001111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100110100";
   IN2_i <= "00001101111011001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110001110";
   IN2_i <= "01010101011101000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110011000";
   IN2_i <= "00010001010111000";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001111110";
   IN2_i <= "00000101110100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001000100";
   IN2_i <= "01000111110000010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011010001";
   IN2_i <= "00000011010001001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000101101";
   IN2_i <= "01110111000011001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010010111";
   IN2_i <= "01110001000010100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100010";
   IN2_i <= "01001001010011000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110001";
   IN2_i <= "01111010000100001";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001110000";
   IN2_i <= "01001001111011111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110100101";
   IN2_i <= "01101111000111000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010100010";
   IN2_i <= "01001101111011001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001001110";
   IN2_i <= "01100100101011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011101111";
   IN2_i <= "00101011011100111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001010110";
   IN2_i <= "01000110101011001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011001001111";
   IN2_i <= "00010110010110001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111110010";
   IN2_i <= "01011001010010100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011010011";
   IN2_i <= "00100001111101010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111100000";
   IN2_i <= "00110011101101101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001100101";
   IN2_i <= "00101101010011110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010110";
   IN2_i <= "00101001011101100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011010001110";
   IN2_i <= "00010011111101110";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001001011";
   IN2_i <= "00010100111111010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101100100";
   IN2_i <= "00001101101001011";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001000011";
   IN2_i <= "01000101100000001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101010101";
   IN2_i <= "01101100110001001";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111101000";
   IN2_i <= "01010010111010110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001111101";
   IN2_i <= "01110001000011000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101000111";
   IN2_i <= "01011100000001010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000100011";
   IN2_i <= "01000010101100111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100011110";
   IN2_i <= "00000011111001010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110011111";
   IN2_i <= "00111000011101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111000001";
   IN2_i <= "01000001101010111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100111001";
   IN2_i <= "01111011100011000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100011000";
   IN2_i <= "00110010101111010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010000000";
   IN2_i <= "01010001111110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010011";
   IN2_i <= "01000111001001001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010000111";
   IN2_i <= "01101100110100011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000111011";
   IN2_i <= "00101111100100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100011111";
   IN2_i <= "01111011010101111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110111000";
   IN2_i <= "00010000110001011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001010010";
   IN2_i <= "01110110110010110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110111111";
   IN2_i <= "01000100001111111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111011011";
   IN2_i <= "01010101110011000";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001010000";
   IN2_i <= "01001100000111100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111001";
   IN2_i <= "01011001100010100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011000111";
   IN2_i <= "01111100011101110";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010111000";
   IN2_i <= "01011010001000010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000100111";
   IN2_i <= "00000101111010101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011001101";
   IN2_i <= "00111000100011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101000010";
   IN2_i <= "01101110010010010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011110101";
   IN2_i <= "00001011001100101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010010110";
   IN2_i <= "00010001000011101";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000111000";
   IN2_i <= "01001001001001001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111100011";
   IN2_i <= "01001010011001000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110010";
   IN2_i <= "01100000011111011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111010101";
   IN2_i <= "00011001000111011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001011011";
   IN2_i <= "01100011011001010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000001000";
   IN2_i <= "00111110010100110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010000100";
   IN2_i <= "00000011101010011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000011010";
   IN2_i <= "00110111100111010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100001110";
   IN2_i <= "00101100100011010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100100000";
   IN2_i <= "00111100110001000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000100110";
   IN2_i <= "00111111011011110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000110001";
   IN2_i <= "00010000000110010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100110";
   IN2_i <= "01101011100101010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111001101";
   IN2_i <= "00000000011111101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000010110";
   IN2_i <= "00110100111000010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110101100";
   IN2_i <= "00010110101010101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110111011011";
   IN2_i <= "00110010101011000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101100010";
   IN2_i <= "01000101101100110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001001001";
   IN2_i <= "00001111001110000";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100000110";
   IN2_i <= "00101110001100110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010111010";
   IN2_i <= "00000101001100111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110010";
   IN2_i <= "00111010101010010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000010010";
   IN2_i <= "00010000001001011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110101100011";
   IN2_i <= "00010110111110010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010110";
   IN2_i <= "00110010010100011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011001101";
   IN2_i <= "00101000011101100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000001000";
   IN2_i <= "00000100101111011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111111000";
   IN2_i <= "01111000101100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101001100";
   IN2_i <= "01110010011011110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011100110";
   IN2_i <= "00111001011100100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100000011";
   IN2_i <= "00001110111111111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001100111";
   IN2_i <= "01001001011100010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001100011";
   IN2_i <= "00101100010011000";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100111011";
   IN2_i <= "01110010001111001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000011010";
   IN2_i <= "01101100110000011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010111001";
   IN2_i <= "00011100001010000";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110110111";
   IN2_i <= "00100010010010100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000111001";
   IN2_i <= "00111001011111101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010100011";
   IN2_i <= "00111111000110010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110111111";
   IN2_i <= "01100101010011011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011000101";
   IN2_i <= "00110110110010100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110101011";
   IN2_i <= "00101101110110011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110111110";
   IN2_i <= "01111111100101010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000011110";
   IN2_i <= "01001001111111011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101100100";
   IN2_i <= "01110010110010000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010011100";
   IN2_i <= "01111000101000100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100000000";
   IN2_i <= "01000010111110100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111111100";
   IN2_i <= "00101101010001010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000011101";
   IN2_i <= "00010110000110101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010011011";
   IN2_i <= "01001011010001101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110010110";
   IN2_i <= "01110110001110000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100011";
   IN2_i <= "00101101001000110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000001011";
   IN2_i <= "01100011110001101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110110101";
   IN2_i <= "01101111011110101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001001001";
   IN2_i <= "00000100101111111";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101010011";
   IN2_i <= "01100011001101100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110011101";
   IN2_i <= "00100101110100111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011101100";
   IN2_i <= "00001111011011000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101011011";
   IN2_i <= "01011101011000100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000001010";
   IN2_i <= "00100001101001001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110011";
   IN2_i <= "00111100111000011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010101101";
   IN2_i <= "00100001110100100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111100011";
   IN2_i <= "01111001010010001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111101010";
   IN2_i <= "01111110000000001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111010111";
   IN2_i <= "01010100010100010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101100101";
   IN2_i <= "01010011001110100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000010111100";
   IN2_i <= "01111100100001101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001100001";
   IN2_i <= "00110100111011000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000111110";
   IN2_i <= "00111101011101110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101110010";
   IN2_i <= "00101110111101010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100011110";
   IN2_i <= "00001011001111000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111111101";
   IN2_i <= "01111001000001101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000101101";
   IN2_i <= "00101100011101110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010111";
   IN2_i <= "00011010000101010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001101111";
   IN2_i <= "00010101110110011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110101110";
   IN2_i <= "00110000011000011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100010111";
   IN2_i <= "01101100100111000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101011011111";
   IN2_i <= "00000101100111010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111111000";
   IN2_i <= "01100100010001101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101101001";
   IN2_i <= "01100000010011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111010110";
   IN2_i <= "00100010111100100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001100001";
   IN2_i <= "00111100000100111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100011111";
   IN2_i <= "00110101100110110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111111011";
   IN2_i <= "00100100001111010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011100110";
   IN2_i <= "00100100110010111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000101101";
   IN2_i <= "01100111001000011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110100110";
   IN2_i <= "01100101100110111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000000010";
   IN2_i <= "00100110100101110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100100";
   IN2_i <= "00111100000100110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010011110";
   IN2_i <= "00000101001100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010110100";
   IN2_i <= "01110110100000110";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110010001";
   IN2_i <= "01100111110011001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010111101";
   IN2_i <= "00001001011101000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100011100";
   IN2_i <= "01111000111000001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100011011";
   IN2_i <= "00100001000001010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110110100";
   IN2_i <= "01001011100001010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000111011";
   IN2_i <= "00001011111000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101010111";
   IN2_i <= "01100100010000001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011110";
   IN2_i <= "00101111011010110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100000000";
   IN2_i <= "00011101000001101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111001011";
   IN2_i <= "01010010111000101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111100001";
   IN2_i <= "00001000100010011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010100000000";
   IN2_i <= "00101001101001100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011110111";
   IN2_i <= "01001101010100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001010000";
   IN2_i <= "00100111111110100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011111000";
   IN2_i <= "00000100011000011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010011110";
   IN2_i <= "01100100001011011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110000110";
   IN2_i <= "00101011000100010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101001001";
   IN2_i <= "01101111000011100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101100100";
   IN2_i <= "00110111010000110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000011000";
   IN2_i <= "01000000001011100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110000101";
   IN2_i <= "01001010110011011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011100100";
   IN2_i <= "01101100001000100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100010101";
   IN2_i <= "01101011111011011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010111";
   IN2_i <= "00010111100001011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001011000";
   IN2_i <= "01011110100010011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110110000";
   IN2_i <= "00110110011010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001010001";
   IN2_i <= "00111001111110001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001010010";
   IN2_i <= "00001001110111110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001101010";
   IN2_i <= "01010001000110100";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001011001";
   IN2_i <= "01010010011100110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010111";
   IN2_i <= "01011110010101110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011000101";
   IN2_i <= "00011111110001000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001001111";
   IN2_i <= "01100011011010011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111110111";
   IN2_i <= "00001001101110001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000010011";
   IN2_i <= "00010110011011111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010100011";
   IN2_i <= "01000101110101001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110111101";
   IN2_i <= "00011001101100010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110111010";
   IN2_i <= "00110110111010101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101001001";
   IN2_i <= "00001100101111000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110100001";
   IN2_i <= "01000111100000011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011011100";
   IN2_i <= "00100100100110011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010100011";
   IN2_i <= "00001111011001110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010010";
   IN2_i <= "01101110011110110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100100001";
   IN2_i <= "01100011110000111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101101110";
   IN2_i <= "01100001110000001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101100001";
   IN2_i <= "00110011000001011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010100100";
   IN2_i <= "01111111011011110";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101100010";
   IN2_i <= "01010010000100010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100000";
   IN2_i <= "01110011111011001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000011100";
   IN2_i <= "01001010001011111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000101010";
   IN2_i <= "00100101001011111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101111110";
   IN2_i <= "00111100100000101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100111110";
   IN2_i <= "01011001001110001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001000000";
   IN2_i <= "00000001000101111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101011010";
   IN2_i <= "01001011011011101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000011101";
   IN2_i <= "01111101111010011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101100010";
   IN2_i <= "00110101010111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110111000";
   IN2_i <= "00101101011011110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101110011";
   IN2_i <= "01100011111100101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110101100";
   IN2_i <= "01001111001100110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100001100";
   IN2_i <= "00110110001011100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101001001";
   IN2_i <= "00110111001110110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001011101";
   IN2_i <= "00101000001110011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110000101";
   IN2_i <= "00011000111010100";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001100101";
   IN2_i <= "01110100110001101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011000001";
   IN2_i <= "01011101110011011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001001111";
   IN2_i <= "00101111000101111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011000000";
   IN2_i <= "01001010010101100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100100111";
   IN2_i <= "01101111000010100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110110010";
   IN2_i <= "01110110000100100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100000";
   IN2_i <= "01100001011111001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110110010";
   IN2_i <= "00010100110001001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011010000";
   IN2_i <= "01110111011111001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001100101";
   IN2_i <= "00011110111110110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110100011";
   IN2_i <= "00010001100010000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101100010";
   IN2_i <= "01100111111011010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011011100";
   IN2_i <= "00111001100000011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101110101";
   IN2_i <= "01100010100000010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101100100";
   IN2_i <= "00101110110001100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101000110";
   IN2_i <= "01100000000101011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000001";
   IN2_i <= "00111000110101010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010110001";
   IN2_i <= "00001011100100101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111001110";
   IN2_i <= "00000011011111001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010011000";
   IN2_i <= "01001000011101100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111011011";
   IN2_i <= "00000001101000111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101110111";
   IN2_i <= "00100000101110011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100001011";
   IN2_i <= "00011011100111111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110000101";
   IN2_i <= "00000001101110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111110011";
   IN2_i <= "00011110011001100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011111101";
   IN2_i <= "00000101110101001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010001101";
   IN2_i <= "00000111110110000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111101000";
   IN2_i <= "00000001101101110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010111111";
   IN2_i <= "01101001111100100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110101";
   IN2_i <= "00010100111010011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100001101";
   IN2_i <= "00000101001100010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001111111";
   IN2_i <= "01111010110001101";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110010";
   IN2_i <= "01101100100011101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111000111";
   IN2_i <= "01100101011010000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101101011";
   IN2_i <= "01001100010101011";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011000111";
   IN2_i <= "00001010100000000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110000100000";
   IN2_i <= "00100100000111011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101111001";
   IN2_i <= "01000001010001101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011100000";
   IN2_i <= "01011100010100110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000010000";
   IN2_i <= "00010001101001011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111110000";
   IN2_i <= "00111111110000000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010010100";
   IN2_i <= "00101010110000100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011000010";
   IN2_i <= "01011001111000011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111010100";
   IN2_i <= "00110000101000001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101100110";
   IN2_i <= "00111100111110010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111101001011";
   IN2_i <= "01100011101110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001010011";
   IN2_i <= "00101000101010000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011110101";
   IN2_i <= "00010101100010010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011111011";
   IN2_i <= "00110111100110100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000011100";
   IN2_i <= "00101110001101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101111010";
   IN2_i <= "01001100010110000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110110100";
   IN2_i <= "01010110011010000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000000";
   IN2_i <= "01010110100111110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101101110";
   IN2_i <= "00000011100100100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101101110000";
   IN2_i <= "00001000000001001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101000000";
   IN2_i <= "01001110110010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111101111";
   IN2_i <= "01000000110110100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000001101";
   IN2_i <= "01001111101110100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010101101";
   IN2_i <= "01110111001010011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001111110";
   IN2_i <= "00110100100010010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000101";
   IN2_i <= "00110001101010100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100101101";
   IN2_i <= "01110110101111001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101101111";
   IN2_i <= "00001001110101001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001100001";
   IN2_i <= "01101101110110000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001110011";
   IN2_i <= "01100011011110001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110000011";
   IN2_i <= "01110101110010101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101101111001";
   IN2_i <= "01010011010100010";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111110111";
   IN2_i <= "00111010110101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100001010";
   IN2_i <= "01110110100111100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000001001";
   IN2_i <= "00111001011010111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001000000";
   IN2_i <= "00101101101011101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001101001110";
   IN2_i <= "00000100000101101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100100111";
   IN2_i <= "00110011000001010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001000100";
   IN2_i <= "00110110111010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001010110";
   IN2_i <= "00010011100000111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101111000";
   IN2_i <= "00001100111110100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000110001";
   IN2_i <= "01111011110100000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100010100110";
   IN2_i <= "00110100010100000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111001011";
   IN2_i <= "00101011000101000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111111001";
   IN2_i <= "00100011000110100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111110110";
   IN2_i <= "01001000001110011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011110000";
   IN2_i <= "01100110001100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100101100";
   IN2_i <= "00011011110100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001111110";
   IN2_i <= "01100011101011000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110100001";
   IN2_i <= "01010010101000001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011011010";
   IN2_i <= "00110111100100111";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000011110";
   IN2_i <= "01011001110110110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111101001";
   IN2_i <= "00011010101010001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111110011";
   IN2_i <= "01000011101111101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000110010";
   IN2_i <= "01011100011000011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000010000";
   IN2_i <= "00110001110001101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010011011";
   IN2_i <= "01000100100100100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110110";
   IN2_i <= "00010110011010001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011001010";
   IN2_i <= "00011110101100010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000110110";
   IN2_i <= "00111111000000010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010101011";
   IN2_i <= "01100010010111110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111100010";
   IN2_i <= "00001110101110000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011110101";
   IN2_i <= "01101101011111011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011011101";
   IN2_i <= "01010101000000010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111011000";
   IN2_i <= "00100100011111000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011000001";
   IN2_i <= "01010010111101100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001000101";
   IN2_i <= "01111100111111111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001011100";
   IN2_i <= "00001000101101011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000000011";
   IN2_i <= "01000001111111101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000111110";
   IN2_i <= "00110101110100101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101100100";
   IN2_i <= "00010011010101010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011000001";
   IN2_i <= "01000111101101110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110010000";
   IN2_i <= "00001100010100001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001001101";
   IN2_i <= "00100111111000000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101100111";
   IN2_i <= "00100100011001101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111001001";
   IN2_i <= "00110011100010110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110101011110";
   IN2_i <= "01001110110010111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001010101";
   IN2_i <= "01100001010010111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010111110";
   IN2_i <= "01111001101110111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010011";
   IN2_i <= "01100110000011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111111011";
   IN2_i <= "01001111110010010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011001111";
   IN2_i <= "01001111010010110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101000101";
   IN2_i <= "01010111100000001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110010011";
   IN2_i <= "01001000100101010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011100000";
   IN2_i <= "01111011101111000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111011111";
   IN2_i <= "00001100100101111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011101001";
   IN2_i <= "01000101101010100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111000000";
   IN2_i <= "00110100000011111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010100110";
   IN2_i <= "00011011101000001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010100111";
   IN2_i <= "00101100001011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000011111";
   IN2_i <= "01111000001101001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010111110";
   IN2_i <= "00001001000101101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110101101";
   IN2_i <= "01100000100011000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100010010";
   IN2_i <= "01000101100000100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110101011";
   IN2_i <= "00110001111011111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101111";
   IN2_i <= "00101001000000010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100110011";
   IN2_i <= "01100000001110111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110101000";
   IN2_i <= "01000000010111100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111110111";
   IN2_i <= "00010001010011110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001001111";
   IN2_i <= "01111100100100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001110000";
   IN2_i <= "00000111001101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011110001";
   IN2_i <= "01100111011011110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110101100";
   IN2_i <= "00101000101010101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001111110";
   IN2_i <= "00101001011010011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001100100";
   IN2_i <= "01001001011001010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011010101";
   IN2_i <= "00110101101000011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100011";
   IN2_i <= "00101110001111101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001011101";
   IN2_i <= "00100010111001011";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100101111";
   IN2_i <= "01000011001010000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101101110";
   IN2_i <= "00101101000011000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110111000";
   IN2_i <= "01110111000100110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110101100";
   IN2_i <= "00011010111101100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011100101";
   IN2_i <= "00110011111001100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111110011";
   IN2_i <= "01111110101100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000010110";
   IN2_i <= "01111010010000101";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000010110";
   IN2_i <= "00010000011011100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010011101";
   IN2_i <= "00010010001010111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011001110";
   IN2_i <= "01010000001101000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010000";
   IN2_i <= "01101010110101011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110010110";
   IN2_i <= "01111000100010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010101101";
   IN2_i <= "01000111110001001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001001000";
   IN2_i <= "00100111011111011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110111000";
   IN2_i <= "01010000111100100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001100111";
   IN2_i <= "01000001110011111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111000011";
   IN2_i <= "01100101101101001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110000011";
   IN2_i <= "00000000010100110";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110011010";
   IN2_i <= "00110001000011110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110111100";
   IN2_i <= "00000000001010110";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110111000";
   IN2_i <= "01011001000001011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000000011";
   IN2_i <= "00111110110110101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111111";
   IN2_i <= "00010001010111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001111011";
   IN2_i <= "00010010111110000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111110001";
   IN2_i <= "01111000001110000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000000110";
   IN2_i <= "01111110001001001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101101";
   IN2_i <= "00001101100011100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110001101";
   IN2_i <= "01100100011100111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001001001";
   IN2_i <= "00011110101001011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110010101";
   IN2_i <= "00110100010001010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110001001";
   IN2_i <= "01100001100111010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010011011";
   IN2_i <= "00100000010010111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011010100";
   IN2_i <= "01001100011010100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111100001";
   IN2_i <= "00101001011100100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101111010";
   IN2_i <= "01010000011110000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010000111";
   IN2_i <= "00110001100100001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100011010101";
   IN2_i <= "01010010101011001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011110001";
   IN2_i <= "00011011111010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010101111";
   IN2_i <= "00111000101011011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101011001";
   IN2_i <= "01111000000110011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000110010";
   IN2_i <= "00001011000110000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001001";
   IN2_i <= "00010011001001011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110110110";
   IN2_i <= "01111111001111101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110110000";
   IN2_i <= "00000011011100010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011100101";
   IN2_i <= "00111010000100111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011100110101";
   IN2_i <= "01011001011100101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000010010";
   IN2_i <= "00100101010010000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111011101";
   IN2_i <= "01101111011100011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110011010";
   IN2_i <= "00111010100101010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011000011";
   IN2_i <= "01001000100000110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110100111";
   IN2_i <= "01011100111011110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011000000";
   IN2_i <= "00111101000100101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001010010";
   IN2_i <= "00010111011000111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101111";
   IN2_i <= "00110110011001100";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111000101";
   IN2_i <= "00111011111010011";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000010000";
   IN2_i <= "01100111111011010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010010011";
   IN2_i <= "01100010111101101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010011111";
   IN2_i <= "00100011011100110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010100111";
   IN2_i <= "00010100001000001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110010110";
   IN2_i <= "01001011101001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011100101";
   IN2_i <= "01100100100011000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011100010";
   IN2_i <= "01111110110000101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011010100";
   IN2_i <= "01101101111100001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000000011";
   IN2_i <= "00001000001001000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100010011";
   IN2_i <= "00101001110010011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011001101";
   IN2_i <= "00110101100111001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010010000";
   IN2_i <= "01000111111001010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011110001";
   IN2_i <= "00010001010110010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011100111";
   IN2_i <= "00110110011101101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100000111";
   IN2_i <= "00010100011101010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110111011";
   IN2_i <= "00110110010011110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111111100";
   IN2_i <= "01000010101011010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111100000";
   IN2_i <= "00010110001010111";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011100100";
   IN2_i <= "01100111111001111";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111011111";
   IN2_i <= "01101111011100000";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010001100";
   IN2_i <= "00110010001110101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111010001";
   IN2_i <= "01111111101010111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111110100";
   IN2_i <= "00001101111011001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000001";
   IN2_i <= "00110010111010111";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111101111111";
   IN2_i <= "01010110001001101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010110110010";
   IN2_i <= "01000001000010111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101110111";
   IN2_i <= "00101100110110101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011100011";
   IN2_i <= "01111001000010110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000011";
   IN2_i <= "01011111101101110";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110011000";
   IN2_i <= "01111001011111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000101110";
   IN2_i <= "01000101101001000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111011111";
   IN2_i <= "00001101011010100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001011101";
   IN2_i <= "01101000011000010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011100011";
   IN2_i <= "01001010111100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011010001";
   IN2_i <= "00110000011011111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011000111";
   IN2_i <= "01101110000101100";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000001111";
   IN2_i <= "00001011110100011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011000";
   IN2_i <= "01101110011101100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011011101";
   IN2_i <= "01011100101111110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010010100";
   IN2_i <= "01100101000001001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110001000";
   IN2_i <= "01010011001011111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101001100";
   IN2_i <= "00100011111011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000111111";
   IN2_i <= "00011000011001000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001001111";
   IN2_i <= "00111100110010111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100110011";
   IN2_i <= "01000011010101111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111001000";
   IN2_i <= "00110000001111001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100111110";
   IN2_i <= "01111110100010101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010010000";
   IN2_i <= "00101111100011111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011000000";
   IN2_i <= "00011011100110111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110110110";
   IN2_i <= "00000010000100011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000001001";
   IN2_i <= "01101001100101000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001100110";
   IN2_i <= "01000110000110111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111101000";
   IN2_i <= "01001110100011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000011010";
   IN2_i <= "00101100011101110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101011110";
   IN2_i <= "00010101100111011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101111100";
   IN2_i <= "01110010010111111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011110011";
   IN2_i <= "00011111011010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101011011";
   IN2_i <= "01011111011001000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111110111";
   IN2_i <= "01110010110000001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101101100";
   IN2_i <= "01001110001001101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010110";
   IN2_i <= "01000100100001000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010110100";
   IN2_i <= "01011010101001000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100010011";
   IN2_i <= "00000011101001000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011111111";
   IN2_i <= "00001001010011000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111011101";
   IN2_i <= "01110110110111000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001010000";
   IN2_i <= "01100001110100110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100000000";
   IN2_i <= "00001010011110100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110011011";
   IN2_i <= "00110010001110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000000001";
   IN2_i <= "00101010001000001";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101010010";
   IN2_i <= "00101100111111011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110111111";
   IN2_i <= "00110101011100111";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000101010";
   IN2_i <= "00010001110111000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001101001";
   IN2_i <= "00001010111110010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011011010";
   IN2_i <= "00111001001011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010100";
   IN2_i <= "00001110111111111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000101000";
   IN2_i <= "00100010100100011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010000110";
   IN2_i <= "00010111010101011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011011000";
   IN2_i <= "00111001011011100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101110110";
   IN2_i <= "01001010100010111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011111111010";
   IN2_i <= "01100101101101110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000000011";
   IN2_i <= "00101010100010111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101010101";
   IN2_i <= "00010001111101000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001110011";
   IN2_i <= "00000110110111000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010100000";
   IN2_i <= "01101111111110011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011001010";
   IN2_i <= "01101111100001111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100000111";
   IN2_i <= "00011100001111000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100010011";
   IN2_i <= "01111010000010000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101110110110";
   IN2_i <= "01110000001100111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011011011";
   IN2_i <= "01011001100101101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011000";
   IN2_i <= "01010000011001011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000001000011";
   IN2_i <= "00110111011011000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100011111";
   IN2_i <= "00110100100000011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000111100";
   IN2_i <= "01000101011011000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110001110";
   IN2_i <= "01100111011010100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011111001";
   IN2_i <= "00011000101000111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010010010";
   IN2_i <= "00000001110011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000100011";
   IN2_i <= "00111001111111011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100101011011";
   IN2_i <= "01101011000101110";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001110010010";
   IN2_i <= "01011011111001000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001001100";
   IN2_i <= "00110010010011100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011001110";
   IN2_i <= "01100011110111001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100010001";
   IN2_i <= "01010110110100011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010111101";
   IN2_i <= "01010110000011110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011110010";
   IN2_i <= "00001110000111000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000101101";
   IN2_i <= "00111001011010001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001011001";
   IN2_i <= "00110011111100001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000000011";
   IN2_i <= "01100011110011011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101001111";
   IN2_i <= "01111100111010101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100110011";
   IN2_i <= "01110110110000001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100000111110";
   IN2_i <= "01001100111111010";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011101111";
   IN2_i <= "01101101110111001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000011010100";
   IN2_i <= "01100001110001011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111001010";
   IN2_i <= "01111100101111101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111100111";
   IN2_i <= "00011001110001100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101111010";
   IN2_i <= "00000000110010101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011010111";
   IN2_i <= "00100110100101010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011101101";
   IN2_i <= "01110010110001001";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000111010";
   IN2_i <= "00001001111010001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100110001";
   IN2_i <= "00110100010000001";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011110001";
   IN2_i <= "01010000000100010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110001";
   IN2_i <= "01100111111110101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110100001";
   IN2_i <= "01101000111010101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101001101";
   IN2_i <= "00010110101100011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110011010";
   IN2_i <= "00110000011110000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000001100";
   IN2_i <= "01110111011011001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110110110";
   IN2_i <= "01000101010011100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001101101101";
   IN2_i <= "00000000100100010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111110111";
   IN2_i <= "01111010111011111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111100110";
   IN2_i <= "00111101101100111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111010101101";
   IN2_i <= "00111011100010011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101001110";
   IN2_i <= "00000000101100101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011100110";
   IN2_i <= "00100001111001001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101010111";
   IN2_i <= "00111111100001111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010100000011";
   IN2_i <= "00001110100101000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111001011";
   IN2_i <= "01011001011111000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111100100";
   IN2_i <= "01101011100111101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010000011";
   IN2_i <= "01000011110001001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010000111";
   IN2_i <= "01010010100001110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100011111";
   IN2_i <= "01010101101000010";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101100101";
   IN2_i <= "01001001111011100";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011001";
   IN2_i <= "00101111000111101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100001010";
   IN2_i <= "00100101000101111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001000111";
   IN2_i <= "01111100100110100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101001110";
   IN2_i <= "01001010101011101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101110011";
   IN2_i <= "01100000001110111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110000001";
   IN2_i <= "01100100001001100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011001101";
   IN2_i <= "00000011011001110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101110111";
   IN2_i <= "00111000001111000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110010101";
   IN2_i <= "00001111000101101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110000100";
   IN2_i <= "00101000011110000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111011110";
   IN2_i <= "00100000100100101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111111100011";
   IN2_i <= "00111001101001000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000011010";
   IN2_i <= "00100100001100111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011100100";
   IN2_i <= "01110111101110110";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101100111";
   IN2_i <= "00101011011100100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101000";
   IN2_i <= "01011001110010110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100111111";
   IN2_i <= "01001101100111111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000100101";
   IN2_i <= "01111110011010100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110011111";
   IN2_i <= "00001111101000100";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010000101";
   IN2_i <= "00010000011100001";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111010100";
   IN2_i <= "01000011110111000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011101000";
   IN2_i <= "00100100011000100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101011000";
   IN2_i <= "01111000010101100";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111110101";
   IN2_i <= "00110100110000001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001011";
   IN2_i <= "00001101011111001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010110101";
   IN2_i <= "01001111101101011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010111101";
   IN2_i <= "01010000101111010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101111010100";
   IN2_i <= "01101100100100100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110010000";
   IN2_i <= "00111010010111011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110001";
   IN2_i <= "00001000011011001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001011";
   IN2_i <= "00100110000110001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001101001";
   IN2_i <= "00011101011001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111110010";
   IN2_i <= "01000100001001000";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100010100";
   IN2_i <= "01100011000111000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111011011";
   IN2_i <= "00101010100101110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000110111";
   IN2_i <= "00001110011110011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011011";
   IN2_i <= "01011000011010010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111000011";
   IN2_i <= "00010000001010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100100000";
   IN2_i <= "01101101000000000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110001100";
   IN2_i <= "00110101111011001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000101001";
   IN2_i <= "01000000011110010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010110";
   IN2_i <= "01111001000010010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100110000";
   IN2_i <= "01101100010001011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110001011";
   IN2_i <= "01011100010101110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101111110";
   IN2_i <= "00000001010011011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111100010";
   IN2_i <= "01011000011100111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100100000";
   IN2_i <= "00001010101100001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100010101";
   IN2_i <= "01001001010110101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001101001";
   IN2_i <= "01000110010001111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010001111";
   IN2_i <= "00110111101001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101101011";
   IN2_i <= "00000100011000111";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101100100";
   IN2_i <= "00100010000001111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111001011";
   IN2_i <= "01101100110001100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001111100";
   IN2_i <= "00011101011100011";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101110010";
   IN2_i <= "01111000011010100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101100111110";
   IN2_i <= "01110100110001000";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000100111";
   IN2_i <= "00011100000001110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111011000000";
   IN2_i <= "00010101011000001";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011010001";
   IN2_i <= "01110011111011011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100001000";
   IN2_i <= "01011111110101111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100101010";
   IN2_i <= "00011111001101100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001100100110";
   IN2_i <= "01001010101110101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001000100";
   IN2_i <= "00001011011100011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110101001";
   IN2_i <= "00100011010111111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010110010";
   IN2_i <= "00010110000011010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011010110";
   IN2_i <= "00101110000010100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110000100";
   IN2_i <= "00011000010011111";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111111111";
   IN2_i <= "00010011110110011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111000011111";
   IN2_i <= "00011110011011010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011011111";
   IN2_i <= "01110100001101111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110000100";
   IN2_i <= "00101001001100110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100010110";
   IN2_i <= "00000101111111011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101011000";
   IN2_i <= "01101000000110101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110010100";
   IN2_i <= "01011001110111110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000111111";
   IN2_i <= "01111110001111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111010001";
   IN2_i <= "01110001111010111";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011100111";
   IN2_i <= "01111110010011100";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110100111";
   IN2_i <= "00111110100011101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010101100";
   IN2_i <= "01101100000101001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011111111111";
   IN2_i <= "01100000100010111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010000000";
   IN2_i <= "00101110111111100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011011011";
   IN2_i <= "01000101010000000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000110111";
   IN2_i <= "01010010111100010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011001101";
   IN2_i <= "01111000100001100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100001110";
   IN2_i <= "01000101111000111";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000000100";
   IN2_i <= "00101100111010000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100110100";
   IN2_i <= "00111110010010010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010110110";
   IN2_i <= "00011110101000111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101111100";
   IN2_i <= "00110111100011100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101011110";
   IN2_i <= "01010110001101101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100001111";
   IN2_i <= "01010110111000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100011000";
   IN2_i <= "01101000110101011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111010110100";
   IN2_i <= "01000110001110111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111101101";
   IN2_i <= "01100100100101010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101110";
   IN2_i <= "01100010011111010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011101101";
   IN2_i <= "01111110100000000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000001000";
   IN2_i <= "01100011000010111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011011111";
   IN2_i <= "00111001100001111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010010100";
   IN2_i <= "00111101000111111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011101111";
   IN2_i <= "00010000000001110";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011010010";
   IN2_i <= "00100101011101101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001110100";
   IN2_i <= "00100110010000110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101001";
   IN2_i <= "00110000000011001";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110101111";
   IN2_i <= "01011010010111111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100111";
   IN2_i <= "01000001101000111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100011111";
   IN2_i <= "01011011000001101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001011010";
   IN2_i <= "01100100110101111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111010011";
   IN2_i <= "00001100000001011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000000000";
   IN2_i <= "00101000011001111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010000111";
   IN2_i <= "00001010000111101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011000001";
   IN2_i <= "00101100000001101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100100011";
   IN2_i <= "00111111011101111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001010011";
   IN2_i <= "01010001001010111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100000000";
   IN2_i <= "00010001100011011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001010101";
   IN2_i <= "00000100100101100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101111001";
   IN2_i <= "01010101000101000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000110001";
   IN2_i <= "01001111011000100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011110000";
   IN2_i <= "01101110010001001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100100101";
   IN2_i <= "01000001101001011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110001101";
   IN2_i <= "01010010000001011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011011101";
   IN2_i <= "00100010011011011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001000011";
   IN2_i <= "00101111000100101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000001011";
   IN2_i <= "01000111011110000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101010000";
   IN2_i <= "00001101100110010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100001001";
   IN2_i <= "00010010101011010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100000100001";
   IN2_i <= "00010001100001000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110011110";
   IN2_i <= "01001010010101111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000100101";
   IN2_i <= "01111000110010011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110101000";
   IN2_i <= "01101001100100111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110010001";
   IN2_i <= "00100111101011100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001001111";
   IN2_i <= "00101101011010110";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111010110";
   IN2_i <= "00000011111010111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111110001";
   IN2_i <= "01011011101010010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010110110";
   IN2_i <= "01001010000011110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010100000";
   IN2_i <= "01010001101101101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010111011001";
   IN2_i <= "01110111010101011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101010100";
   IN2_i <= "01010111001011001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101111101";
   IN2_i <= "01001100010100011";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010001001";
   IN2_i <= "01110111011111001";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101011111";
   IN2_i <= "00001100001011011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011010";
   IN2_i <= "00000111000101100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101011111100";
   IN2_i <= "00100000011101110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000010000";
   IN2_i <= "01000111011110001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101101011100";
   IN2_i <= "00100101110001001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011010111";
   IN2_i <= "01011010101000000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111101110";
   IN2_i <= "01101000101101001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001100100";
   IN2_i <= "00111011100111110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111001000111";
   IN2_i <= "01001011101101101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111010110010";
   IN2_i <= "01110101000101000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011100011";
   IN2_i <= "01110011011001100";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000011111000";
   IN2_i <= "00111001101010001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000001000";
   IN2_i <= "01100011101001101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100101001";
   IN2_i <= "00101100100101000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110011101";
   IN2_i <= "01110001111011110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010000000110";
   IN2_i <= "00111111011010010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111100000";
   IN2_i <= "00011010101001111";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111000111111";
   IN2_i <= "00110010011010111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101001100";
   IN2_i <= "01111010110011001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001011011";
   IN2_i <= "01101101001001110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011111001";
   IN2_i <= "00111100001000101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110110";
   IN2_i <= "00011111110101111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001110000";
   IN2_i <= "01100001010011000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010101101";
   IN2_i <= "00010010011001010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010101101";
   IN2_i <= "01001111101011001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101000111";
   IN2_i <= "00100001100011000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111010";
   IN2_i <= "01111101101101011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111001000";
   IN2_i <= "00000100100000101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110101100";
   IN2_i <= "00011000001111011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000001111";
   IN2_i <= "01111110001010100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111010001";
   IN2_i <= "00110100110100001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000010110";
   IN2_i <= "01110111001101000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000110";
   IN2_i <= "01111000001101011";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000000000";
   IN2_i <= "01101001101101100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011101111";
   IN2_i <= "00011000010111100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100011";
   IN2_i <= "00001010011101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111100000100";
   IN2_i <= "01011010101100000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110110001";
   IN2_i <= "01011001101110001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011001011";
   IN2_i <= "00110001110010110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001111110";
   IN2_i <= "01101110111111010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010110101";
   IN2_i <= "00101000101101110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100100011";
   IN2_i <= "01101001000010101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000101110";
   IN2_i <= "00111001100110001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111110110001";
   IN2_i <= "01010101100000100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111011101";
   IN2_i <= "00001111110101100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101111010";
   IN2_i <= "01111100101110100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010100000";
   IN2_i <= "01111000100001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101111100111";
   IN2_i <= "01010111000001010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000000010";
   IN2_i <= "00011110010001110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100100011";
   IN2_i <= "01000100100011101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101011001";
   IN2_i <= "01111010011001011";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101001101";
   IN2_i <= "00100101000111001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001010100";
   IN2_i <= "00110110110110011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011110011010";
   IN2_i <= "01101101000101100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001001010";
   IN2_i <= "00111010011000111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110100111";
   IN2_i <= "00010101110101111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010111100110";
   IN2_i <= "01111110100001010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110001000";
   IN2_i <= "01101111000100101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110000";
   IN2_i <= "00011001011001111";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101101101";
   IN2_i <= "01010011011011011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001000111";
   IN2_i <= "00111011000100100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111000111";
   IN2_i <= "00111010100000010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011010010011";
   IN2_i <= "01000101101101101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010100101";
   IN2_i <= "01110010101000110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011001000";
   IN2_i <= "00101010110010101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110111110";
   IN2_i <= "01100101111101010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011111111011";
   IN2_i <= "00000111010000010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111100000";
   IN2_i <= "00101100101000010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001111001";
   IN2_i <= "00011111011100011";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100100001";
   IN2_i <= "00001101101111001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010101111001";
   IN2_i <= "00001001011010101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010000011";
   IN2_i <= "01000001111011010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110000101";
   IN2_i <= "00001001100100101";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101111011";
   IN2_i <= "01011100011011011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000110000111";
   IN2_i <= "00000110000110111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101101110";
   IN2_i <= "00011010010010100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101101001";
   IN2_i <= "01000110100110110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100000000";
   IN2_i <= "01110000011001011";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000001010";
   IN2_i <= "01010110011110111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110001010";
   IN2_i <= "00101100011001011";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000000000";
   IN2_i <= "00110110110100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011000101";
   IN2_i <= "01110100001111111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100111011";
   IN2_i <= "01000101011011101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110000101";
   IN2_i <= "00110001111011000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010101101";
   IN2_i <= "00001001001111000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010101111";
   IN2_i <= "00100110000000111";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101001010";
   IN2_i <= "00100100001110000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100101010";
   IN2_i <= "00001011010101001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001010010";
   IN2_i <= "01110100110011010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100011110";
   IN2_i <= "01001101001010011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100101011011";
   IN2_i <= "00100001011100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100001110";
   IN2_i <= "01111011111111010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010100001";
   IN2_i <= "01001111100001110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000111001";
   IN2_i <= "01101100110000100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011011111001";
   IN2_i <= "01100111101110011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010000110001";
   IN2_i <= "00111000110010100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101010001";
   IN2_i <= "00011100010100111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100100010";
   IN2_i <= "00000001000001001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111000101";
   IN2_i <= "00101010110101010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111101010";
   IN2_i <= "01000111110010101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100000001";
   IN2_i <= "00010000100010001";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111110101";
   IN2_i <= "01011100001111000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111110001";
   IN2_i <= "00111100001011010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101100001";
   IN2_i <= "01111100000100101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000100101";
   IN2_i <= "01111010010010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110000000";
   IN2_i <= "00110001010111101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111011100";
   IN2_i <= "01111100101000110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111000010110";
   IN2_i <= "00110100101101011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001100101";
   IN2_i <= "01001010000111101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111011011000";
   IN2_i <= "01111100110000010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011110001";
   IN2_i <= "00110111100011010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000010110101";
   IN2_i <= "00011001000110000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110010011";
   IN2_i <= "00110001111101010";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011110001";
   IN2_i <= "00110001101000101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010111";
   IN2_i <= "00010110111001001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100001010";
   IN2_i <= "00101111000111100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100100101";
   IN2_i <= "01100101101010000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101010001";
   IN2_i <= "01110111110010000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010001101011";
   IN2_i <= "00011101100110100";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001010101";
   IN2_i <= "00001011001111101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111000011";
   IN2_i <= "01100001001001111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100010111";
   IN2_i <= "01101101011100000";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011001110";
   IN2_i <= "00011000001011001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111101000";
   IN2_i <= "00000011101111101";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010010001";
   IN2_i <= "01000010111001111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011111110010";
   IN2_i <= "01101101110010110";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111000100";
   IN2_i <= "00101011001100101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101000111";
   IN2_i <= "01100011111101101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010011111";
   IN2_i <= "01000100011100110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011011111";
   IN2_i <= "00110010100100101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111000100001";
   IN2_i <= "00010111100101001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110011001";
   IN2_i <= "01001000011111001";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011011011";
   IN2_i <= "00000011111001101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100100010";
   IN2_i <= "01101111010110001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110100111";
   IN2_i <= "00010100101011000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101000011";
   IN2_i <= "01001001001001010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101001000";
   IN2_i <= "01111001100010001";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000111111";
   IN2_i <= "01110101000111111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100101001";
   IN2_i <= "01101000001111101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111110";
   IN2_i <= "01110001010001100";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001010011";
   IN2_i <= "00011110110010000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000110000";
   IN2_i <= "00010111101000010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000010001";
   IN2_i <= "01010011101011010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110000010";
   IN2_i <= "00110100010010111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111011001";
   IN2_i <= "00010001101010001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111000001110";
   IN2_i <= "01100111110111101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100000110";
   IN2_i <= "00100101100000001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011100110";
   IN2_i <= "00010111010110010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110000000000";
   IN2_i <= "00000111111101001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101110000";
   IN2_i <= "00000001001101000";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001111011101";
   IN2_i <= "00000001010111100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010100101";
   IN2_i <= "01111001000111010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000010001";
   IN2_i <= "00100101111011101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011011000";
   IN2_i <= "01011010001101111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010110110";
   IN2_i <= "00011101010011011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110100000";
   IN2_i <= "00100100101010111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110010111110";
   IN2_i <= "00010101101111111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010011100";
   IN2_i <= "00011000001011011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000000101";
   IN2_i <= "01011011010010110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000101001";
   IN2_i <= "01001110110101100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100010011111";
   IN2_i <= "00011101111101110";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100000100";
   IN2_i <= "01010011001110000";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111001011";
   IN2_i <= "01010111111010000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001000100";
   IN2_i <= "00111010111011000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010101110";
   IN2_i <= "00110010101111011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111010011";
   IN2_i <= "01000001000101010";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111011000";
   IN2_i <= "00010100001111101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001000110";
   IN2_i <= "01010101111100010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101000";
   IN2_i <= "00011100100011011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101010";
   IN2_i <= "00100101011100001";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011001";
   IN2_i <= "00000011110101111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110111010";
   IN2_i <= "01101110011101100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001100111110";
   IN2_i <= "01000010000001100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000011100";
   IN2_i <= "00101010000010011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101110101010";
   IN2_i <= "00100111000010000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001010100";
   IN2_i <= "00010100001111110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110110011";
   IN2_i <= "01001001000100100";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011010001";
   IN2_i <= "01110101110001101";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001010000";
   IN2_i <= "00100010101010000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001100011";
   IN2_i <= "00101100100101111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111001000";
   IN2_i <= "01111000011111011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111100111";
   IN2_i <= "01000001111011110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011111000111";
   IN2_i <= "00010010111000100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011001011101";
   IN2_i <= "00111000000000110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110000110";
   IN2_i <= "00111101111111100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110111001100";
   IN2_i <= "00011001110001111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101110100";
   IN2_i <= "00100110011010101";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110111001";
   IN2_i <= "01010101111001101";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001110000";
   IN2_i <= "01111001110110100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110011111100";
   IN2_i <= "00011111101100111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001000001001";
   IN2_i <= "00010110111001010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001010110";
   IN2_i <= "01001000110110010";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110100100000";
   IN2_i <= "00001111011100001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110101000";
   IN2_i <= "00110101110100001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011010111";
   IN2_i <= "00000010010000011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011011010";
   IN2_i <= "00010000011100101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101001010";
   IN2_i <= "01010000000111100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011001001";
   IN2_i <= "01001000111100011";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001110011";
   IN2_i <= "01110000011111100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001110110";
   IN2_i <= "00011110000011110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010001100";
   IN2_i <= "01110000110011010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011000100";
   IN2_i <= "01101110101110001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010001000010";
   IN2_i <= "01111000111011101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100111010110";
   IN2_i <= "01001100110010101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011000000";
   IN2_i <= "00010000011100110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101011000";
   IN2_i <= "00100000110100010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001111010";
   IN2_i <= "01000001011001100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101100";
   IN2_i <= "01111001000100111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011100010";
   IN2_i <= "00011000001100001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011011010";
   IN2_i <= "01011011001000010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001100011";
   IN2_i <= "00100101001100100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010111101";
   IN2_i <= "00001000000000101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110110100100";
   IN2_i <= "00010011100111010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111000111";
   IN2_i <= "00001100101000001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111111";
   IN2_i <= "01011010000010011";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100010111";
   IN2_i <= "00010110000000110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000100100";
   IN2_i <= "00011101011011101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100111";
   IN2_i <= "01100011001010000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010001001";
   IN2_i <= "00111110000000100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100000100";
   IN2_i <= "00011111100100110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011011";
   IN2_i <= "00001110001010010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010000000";
   IN2_i <= "01111101100111101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110101";
   IN2_i <= "00000111111110011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011011000";
   IN2_i <= "00110111000010011";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111101101";
   IN2_i <= "01010001000110101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100001011";
   IN2_i <= "00110011010000101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100101111";
   IN2_i <= "01011000101001000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010000000";
   IN2_i <= "01000100110100110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001110111000";
   IN2_i <= "00001001101110001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010011010001";
   IN2_i <= "01001001110101111";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011100010";
   IN2_i <= "00111011101011011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010000101";
   IN2_i <= "00110000100101100";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001111111";
   IN2_i <= "01101111010100101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111001110";
   IN2_i <= "00000001111001110";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100000110";
   IN2_i <= "00011111011111000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010100011";
   IN2_i <= "00101010101111001";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111010101";
   IN2_i <= "01001100110111100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100111011";
   IN2_i <= "00100000011000100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110110000";
   IN2_i <= "01010100011111001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111110100";
   IN2_i <= "01101010101111010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001100010";
   IN2_i <= "01101101100100001";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111110101100";
   IN2_i <= "00101111010111000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001000010";
   IN2_i <= "01100100001010010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100000010";
   IN2_i <= "01111001100110011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011001001110";
   IN2_i <= "01001001110111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000011001";
   IN2_i <= "00111110010000001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011111011";
   IN2_i <= "01110010010000011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000110100001";
   IN2_i <= "00110010011101001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011101001";
   IN2_i <= "01100000111111010";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010000100";
   IN2_i <= "01110000101110011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101011111";
   IN2_i <= "00110101100010111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100110111";
   IN2_i <= "00101010010101111";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011000101";
   IN2_i <= "00011100101111001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001000101";
   IN2_i <= "00011110101001110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010010111";
   IN2_i <= "00111111001100101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101100001010";
   IN2_i <= "00000010110100010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110101000";
   IN2_i <= "00000110111000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101111111";
   IN2_i <= "01100010100101111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000000001";
   IN2_i <= "00101100111101001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101111010100";
   IN2_i <= "01000001010000000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010000111";
   IN2_i <= "01110101100101110";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111100111";
   IN2_i <= "01111111100110101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010001101";
   IN2_i <= "01001110000001101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001101001";
   IN2_i <= "00000101100110001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101001010110";
   IN2_i <= "01001111000100101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101001101001";
   IN2_i <= "00111001011100101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011110100110";
   IN2_i <= "00111010101111100";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111000000";
   IN2_i <= "01110000101000110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110110100";
   IN2_i <= "01000000010000000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010100011";
   IN2_i <= "01111001000011011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000100101";
   IN2_i <= "01010011101110101";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000000110";
   IN2_i <= "00111000111101000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110111111";
   IN2_i <= "01000110010010000";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101100000";
   IN2_i <= "01111001001110110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010011111000";
   IN2_i <= "00111010110000111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001001";
   IN2_i <= "00001101010100101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011011010";
   IN2_i <= "01111011101011101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111011101111";
   IN2_i <= "01011001100011011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101010111111";
   IN2_i <= "00111011010100000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010100010";
   IN2_i <= "00101011101111010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101110000";
   IN2_i <= "00011011010101101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001111110";
   IN2_i <= "00101011111100000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111001001100";
   IN2_i <= "01001100001010010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010101001";
   IN2_i <= "01100111110000110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010100110";
   IN2_i <= "01111001011010111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100101011000";
   IN2_i <= "01101010011111101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001010111";
   IN2_i <= "01101011110001110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011000110101";
   IN2_i <= "01100000001100100";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001110101";
   IN2_i <= "01000100110010101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000000110";
   IN2_i <= "01100101001001110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101110";
   IN2_i <= "00111001010101011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010000011010";
   IN2_i <= "01001100110101011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101000010";
   IN2_i <= "00101010011001001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011101110110";
   IN2_i <= "00011100110001000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111010100";
   IN2_i <= "01011001100011010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011101100";
   IN2_i <= "00000011001001101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111001111";
   IN2_i <= "00101010110100101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110001011";
   IN2_i <= "00010111010101101";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001000100";
   IN2_i <= "00011111111101010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000011001";
   IN2_i <= "01111011111101001";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111001000";
   IN2_i <= "00000111101010101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110110010";
   IN2_i <= "01000010010001000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101011111010";
   IN2_i <= "01001010011011000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111101000101";
   IN2_i <= "01100100000001110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101110000011";
   IN2_i <= "00000010001010001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010010011";
   IN2_i <= "01111011011100011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100010011101";
   IN2_i <= "00000011110011101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010101101";
   IN2_i <= "01111111011100000";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000010100111";
   IN2_i <= "01110101101000111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101100110";
   IN2_i <= "01000111001101101";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100011010";
   IN2_i <= "01111100101110010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100010111";
   IN2_i <= "01101100010001100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101100101";
   IN2_i <= "00000110100111111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111010001";
   IN2_i <= "01010010000001110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111001101";
   IN2_i <= "00000101100001011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011111010";
   IN2_i <= "01100101110100010";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000110011";
   IN2_i <= "01011101010111000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111110011101";
   IN2_i <= "00101110010100101";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101111101";
   IN2_i <= "01101100100010011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010010000";
   IN2_i <= "01001100110110010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001000010000";
   IN2_i <= "00110111110110100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011111000";
   IN2_i <= "01100100100111110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001101111001";
   IN2_i <= "01101110110110001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110010110";
   IN2_i <= "01100000100010110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111110101";
   IN2_i <= "00111010011101101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010110101";
   IN2_i <= "01110111001110001";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100000101001";
   IN2_i <= "01100011110010101";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100001010";
   IN2_i <= "00110011101000000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100110101";
   IN2_i <= "00011110110001011";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100011";
   IN2_i <= "00011010001001010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000010101";
   IN2_i <= "01000001011101011";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001010000";
   IN2_i <= "01010011010001011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000111011";
   IN2_i <= "01011100110011100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111110010";
   IN2_i <= "00111000000010110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110101101";
   IN2_i <= "00001010100000111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010011010";
   IN2_i <= "00010010101100100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111111111";
   IN2_i <= "01000010011101101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011101000";
   IN2_i <= "01010101111000001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000000011";
   IN2_i <= "01110001001110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111101011";
   IN2_i <= "00010101001100100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011000010";
   IN2_i <= "01111001101000010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100111010000";
   IN2_i <= "00001101000001011";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000101100";
   IN2_i <= "00011110000111110";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100001101";
   IN2_i <= "01111000110010100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011101000001";
   IN2_i <= "01010001000100110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111101010";
   IN2_i <= "00001011101110000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110111011";
   IN2_i <= "01000000110111110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100001011";
   IN2_i <= "00011001001001111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110111010";
   IN2_i <= "00011000000011011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001100001";
   IN2_i <= "01101100011101000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101001000";
   IN2_i <= "01010100000001000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000000000010";
   IN2_i <= "00010111000110111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110000111";
   IN2_i <= "01100100000010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010110011111";
   IN2_i <= "00100100110001000";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010010100";
   IN2_i <= "00010101000010000";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010011010";
   IN2_i <= "01101110000101000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111011100100";
   IN2_i <= "00001000101010000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111000000";
   IN2_i <= "01010111010001111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111011010";
   IN2_i <= "00001111100010010";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011100010";
   IN2_i <= "00001111110011000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110100000";
   IN2_i <= "00010011011010111";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000100101";
   IN2_i <= "00101101101111010";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100101110";
   IN2_i <= "00111011110101001";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100010011";
   IN2_i <= "00111011001100110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000001000";
   IN2_i <= "00100100110011001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111000101";
   IN2_i <= "00110111111010111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001011101";
   IN2_i <= "00010000001100111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100001111";
   IN2_i <= "00111100001111001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010011111100";
   IN2_i <= "00011110010110011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010011101";
   IN2_i <= "01001100110000011";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100010101";
   IN2_i <= "01001100110011110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100010110";
   IN2_i <= "00101100001101110";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101001001";
   IN2_i <= "00101010111000100";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010111011010";
   IN2_i <= "00011001011100101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100001100111";
   IN2_i <= "01011101000000011";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011110110";
   IN2_i <= "00010110011011111";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010100110";
   IN2_i <= "01110100100000000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001111001";
   IN2_i <= "00100001010010000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000001001";
   IN2_i <= "01101101100011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000010101";
   IN2_i <= "01100100011110110";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110010101";
   IN2_i <= "01101001000010110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001000111";
   IN2_i <= "01000001111011100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010001111";
   IN2_i <= "00001000101000010";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010100111";
   IN2_i <= "00000000010011010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101010110";
   IN2_i <= "00101110110101000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010110010110";
   IN2_i <= "00111010110111000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110101111";
   IN2_i <= "00100010111100011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011111100";
   IN2_i <= "00000111000101010";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011101101011";
   IN2_i <= "00011001111110110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110011100";
   IN2_i <= "01000100110001001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001000100";
   IN2_i <= "00001101101011100";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001101001";
   IN2_i <= "00111000011000011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010110111";
   IN2_i <= "00101111011010011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010010111110";
   IN2_i <= "00101000111011110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110111110";
   IN2_i <= "00010011101101001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011111001";
   IN2_i <= "00001010001011001";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000110101";
   IN2_i <= "00110110100011110";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011000000";
   IN2_i <= "00110011000100101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010101100";
   IN2_i <= "00110101111110000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010000010";
   IN2_i <= "01101010011011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001011100";
   IN2_i <= "00110110000111111";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110100010001";
   IN2_i <= "01011101000111011";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110010100";
   IN2_i <= "00000100001101001";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110001011";
   IN2_i <= "01110001101000101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001010010101";
   IN2_i <= "01011111001011010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111010100";
   IN2_i <= "01101011100110010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110010010";
   IN2_i <= "00000101100000110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111011011";
   IN2_i <= "01111010111100110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000101111111";
   IN2_i <= "01101100001111101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100001";
   IN2_i <= "01110000100110101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101101001";
   IN2_i <= "00011110101011101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111100001";
   IN2_i <= "00000011000000010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101001010";
   IN2_i <= "01111000010101001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011111100";
   IN2_i <= "01010010010110101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010000011";
   IN2_i <= "01100111100101111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100111010";
   IN2_i <= "01100010100110001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000111001";
   IN2_i <= "01110011100100000";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110001011001";
   IN2_i <= "01000011100101000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100000100011";
   IN2_i <= "00011101111101011";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011110001101";
   IN2_i <= "01111000011111111";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110101101";
   IN2_i <= "00111100100110001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110011010011";
   IN2_i <= "01101111101100110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111010001";
   IN2_i <= "00110000101000101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110110001";
   IN2_i <= "00100000001101000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101101000";
   IN2_i <= "01001101011001101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110110110101";
   IN2_i <= "01100110100000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001010010";
   IN2_i <= "00001000111101011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010011010";
   IN2_i <= "01000010101111011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011010100";
   IN2_i <= "00101111100000000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101000110";
   IN2_i <= "00100111101010010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010001101";
   IN2_i <= "01110100111000000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100010011";
   IN2_i <= "01100001001110010";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100001101010";
   IN2_i <= "00011010000000000";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001011101";
   IN2_i <= "00000111100100000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001111000010";
   IN2_i <= "01011011110100100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000100011";
   IN2_i <= "01010101010110011";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110101100";
   IN2_i <= "00101101010101001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111010100";
   IN2_i <= "00111010000101010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111111000100";
   IN2_i <= "01011000110000010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110000001";
   IN2_i <= "00011000001110011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100001101";
   IN2_i <= "01100100101000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101100011";
   IN2_i <= "01011110001010101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001101001110";
   IN2_i <= "01111010110011100";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111010101";
   IN2_i <= "01000001011011100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101101111";
   IN2_i <= "00000111111000100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001000010000";
   IN2_i <= "00101011000001100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111100100";
   IN2_i <= "01111110100011110";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101000010";
   IN2_i <= "00000101111101011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001010001";
   IN2_i <= "00100000100011111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111101101";
   IN2_i <= "00001110101011011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000011100101";
   IN2_i <= "00001111111010000";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011010111";
   IN2_i <= "00111101010110011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001000010";
   IN2_i <= "00011110010011110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000111101";
   IN2_i <= "00100101100010110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011110";
   IN2_i <= "00000010110011001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001110110";
   IN2_i <= "00011101101110011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101011110";
   IN2_i <= "01111110001100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000110011";
   IN2_i <= "01011100011111011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000100111";
   IN2_i <= "01001011000110101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000111110";
   IN2_i <= "00101000001110101";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010101111";
   IN2_i <= "00010100011111001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101110100";
   IN2_i <= "01111110101100011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101000110";
   IN2_i <= "00100011010010110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100111110";
   IN2_i <= "00001001011101111";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111101100";
   IN2_i <= "00101010011000001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110000001011";
   IN2_i <= "01110111100100110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001001100100";
   IN2_i <= "01000101011000100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000110010";
   IN2_i <= "01000100000110101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000100000";
   IN2_i <= "00101110010101010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001111010";
   IN2_i <= "01100110111011101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110000111000";
   IN2_i <= "01100011101101101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101010001110";
   IN2_i <= "01010110111010100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110101001";
   IN2_i <= "01011110010010010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101100110001";
   IN2_i <= "01000111101111011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101110001";
   IN2_i <= "01000011111110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001111101100";
   IN2_i <= "00101101000010011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100000000";
   IN2_i <= "00000100010000111";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111000110";
   IN2_i <= "01111100000100011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111011010";
   IN2_i <= "00010111011011110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001011110110";
   IN2_i <= "01101000100001110";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000110011";
   IN2_i <= "00100011111011101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100010000";
   IN2_i <= "00010011011010000";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110001000101";
   IN2_i <= "00100101010001011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111110110";
   IN2_i <= "00011001111110111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101101011";
   IN2_i <= "01110001100111100";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111010010";
   IN2_i <= "00010111100110010";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101110001";
   IN2_i <= "00110001010111001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110011110";
   IN2_i <= "00110000101110000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010110001";
   IN2_i <= "00001110010110110";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000100101";
   IN2_i <= "01011010001101011";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000110000110";
   IN2_i <= "00001001011001101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000101001";
   IN2_i <= "00010000111010111";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100001";
   IN2_i <= "00010000101011101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001001000";
   IN2_i <= "01110001010010111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110010010";
   IN2_i <= "01110111100000011";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000000101";
   IN2_i <= "00010100111000101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011100111";
   IN2_i <= "00010000010001100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001101100";
   IN2_i <= "01011011011010110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101101101";
   IN2_i <= "01000100000110101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011001111111";
   IN2_i <= "00111110000011110";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010110000";
   IN2_i <= "01111111001001110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010101010100";
   IN2_i <= "00000011111100000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000011110001";
   IN2_i <= "01111011010011011";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010100011";
   IN2_i <= "00010101001110101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000010111";
   IN2_i <= "01011111011011111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000101000";
   IN2_i <= "01000000000011000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000001010";
   IN2_i <= "01101000010000001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100000100010";
   IN2_i <= "00011101101100000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001000100";
   IN2_i <= "01100010001000111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010100000";
   IN2_i <= "01111111110001010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010110011";
   IN2_i <= "01001111111000010";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011000000";
   IN2_i <= "00000110110100100";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101100001";
   IN2_i <= "01000110110111110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101000110";
   IN2_i <= "00001101101011000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010010111110";
   IN2_i <= "00010001010011100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001001111010";
   IN2_i <= "00110010000001101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011111110";
   IN2_i <= "00111010001011101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010001000";
   IN2_i <= "00110001011010000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101011001";
   IN2_i <= "01110100101111100";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110110011100";
   IN2_i <= "00111100010010111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011101011000";
   IN2_i <= "00100011000010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011111010";
   IN2_i <= "00000000011011001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111001001";
   IN2_i <= "01001000000101010";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111011001";
   IN2_i <= "01011101011101101";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100100111";
   IN2_i <= "00011110100100111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000101110";
   IN2_i <= "00100001110011101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111100111000";
   IN2_i <= "01111111011011010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111001111001";
   IN2_i <= "00100001011100100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011001001011";
   IN2_i <= "01001100100000011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101100000";
   IN2_i <= "01100111000100111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010110010";
   IN2_i <= "00001111011000000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010101101000";
   IN2_i <= "00000011011001011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101011101";
   IN2_i <= "00011110110100100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011100010010";
   IN2_i <= "00101010010010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100101110";
   IN2_i <= "00110010010100000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110001100";
   IN2_i <= "00111101000010011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011001111";
   IN2_i <= "00101000011110110";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010001010000";
   IN2_i <= "01011110010011001";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000001111000";
   IN2_i <= "01101010010111001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100100100";
   IN2_i <= "01011000110000000";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100011001";
   IN2_i <= "00010010100110110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100001110";
   IN2_i <= "00111101000111111";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101110100011";
   IN2_i <= "00101100101101101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101010001010";
   IN2_i <= "01100101001100100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111010011";
   IN2_i <= "01111110100111010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100100110000";
   IN2_i <= "00111111001111100";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100000111";
   IN2_i <= "01011100101000110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100100101100";
   IN2_i <= "01010001010101111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101101001111";
   IN2_i <= "00111110100001001";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101001010";
   IN2_i <= "01001011111111001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011000000";
   IN2_i <= "01110011111110010";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100110001";
   IN2_i <= "01110000000010011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100001111";
   IN2_i <= "01011100010011100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100000";
   IN2_i <= "01011110100000010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011011011";
   IN2_i <= "00001010000011010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010100100";
   IN2_i <= "01000000110010100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101110001";
   IN2_i <= "01110100010110101";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000101101";
   IN2_i <= "01010001000011100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100100101001";
   IN2_i <= "01101101111100000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000110010111";
   IN2_i <= "00000111010100001";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101101111";
   IN2_i <= "00000101010011000";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100011000010";
   IN2_i <= "00011111011111100";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001110000";
   IN2_i <= "00101100100110010";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101101000";
   IN2_i <= "01100100001000011";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000101100011";
   IN2_i <= "00010011000110001";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010011111";
   IN2_i <= "01000011101100001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100110000011";
   IN2_i <= "01111011010001010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000011";
   IN2_i <= "01011101110110001";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111000000";
   IN2_i <= "00000000000011111";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010011001";
   IN2_i <= "01010001000011100";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011111011000";
   IN2_i <= "01001010001101001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010000010110";
   IN2_i <= "00110010100110010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110101111";
   IN2_i <= "00100111111101101";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000011111";
   IN2_i <= "01010010101011010";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000100010001";
   IN2_i <= "00001110011010010";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101001";
   IN2_i <= "00101000000001001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111100110";
   IN2_i <= "00110111010100101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111001110111";
   IN2_i <= "00001101010101000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001110001";
   IN2_i <= "00110000101010010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101111100110";
   IN2_i <= "00110000101110100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001000011111";
   IN2_i <= "01010100011110001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010011101";
   IN2_i <= "00101000111100100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010001111";
   IN2_i <= "01010101111110001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000111010";
   IN2_i <= "00010010000110001";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101100000";
   IN2_i <= "00111110111100111";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010010010010";
   IN2_i <= "00011100111001010";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101011000101";
   IN2_i <= "01110000110110000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010010010001";
   IN2_i <= "00111101000000111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000000001111";
   IN2_i <= "00100111010000000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101101100";
   IN2_i <= "01000001100011100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000111000111";
   IN2_i <= "00001110110010010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100101011";
   IN2_i <= "01100110001000100";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011000011";
   IN2_i <= "01100011001100011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110010001010";
   IN2_i <= "01001101100111011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011100110101";
   IN2_i <= "01010100001001100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101000111";
   IN2_i <= "01011101010100101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010110101";
   IN2_i <= "01101101100011011";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101111000101";
   IN2_i <= "01111101101111001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111100100101";
   IN2_i <= "01110101010100101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110001001";
   IN2_i <= "00110100100001101";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111100100";
   IN2_i <= "01101100101000001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011111101";
   IN2_i <= "01000110000011110";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100101101001";
   IN2_i <= "00110101000011101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101010001";
   IN2_i <= "00010100101011010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110001001001";
   IN2_i <= "00010101000000001";
   IN3_i <= "0011110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100011001100";
   IN2_i <= "01000010011111010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000010100";
   IN2_i <= "01001100000101010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100100011";
   IN2_i <= "00101111101000011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100011001";
   IN2_i <= "01110001111110001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001111000";
   IN2_i <= "00001010000000110";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000101110";
   IN2_i <= "00011011100100101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111100011";
   IN2_i <= "01000010110101110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111011101001";
   IN2_i <= "00000101110011001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110001010110";
   IN2_i <= "01000010111001101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100100101";
   IN2_i <= "00011111101110100";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010111010";
   IN2_i <= "00100010111101100";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011011111";
   IN2_i <= "00000010000001000";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001101101100";
   IN2_i <= "00001111110111010";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101111011";
   IN2_i <= "01010100110010000";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100000110";
   IN2_i <= "01011111110111100";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101011001";
   IN2_i <= "01010111001000111";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111010011001";
   IN2_i <= "01100101011110110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101111011";
   IN2_i <= "01100111010101000";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010100011";
   IN2_i <= "00101010100101000";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001111000101";
   IN2_i <= "01111110011110000";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000010011";
   IN2_i <= "01001101110000000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010101000001";
   IN2_i <= "01011101001100111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100001101101";
   IN2_i <= "00000000101100111";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100000011";
   IN2_i <= "00101110011111101";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001110011101";
   IN2_i <= "01100110011111110";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000100001110";
   IN2_i <= "01111000011011100";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001000";
   IN2_i <= "00100100100110011";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101000110";
   IN2_i <= "01010011001000111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011011010";
   IN2_i <= "01001101011101010";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010111001";
   IN2_i <= "00101010011000011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001001101110";
   IN2_i <= "00000110000110111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111110110110";
   IN2_i <= "01011011111011110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111100100101";
   IN2_i <= "01000010011111100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001000101";
   IN2_i <= "00010111100111111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110110110";
   IN2_i <= "01100011000111000";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001000111";
   IN2_i <= "00000001001101000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111101111";
   IN2_i <= "00011000000111000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101011100001";
   IN2_i <= "00010011100110011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110011101110";
   IN2_i <= "00100100101110101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110010001";
   IN2_i <= "01101001111011010";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100101010";
   IN2_i <= "01100100111001010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101110101111";
   IN2_i <= "01101011110110000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101001110000";
   IN2_i <= "00101010101110010";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110111010";
   IN2_i <= "00100111100001000";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000110001";
   IN2_i <= "00110101100001111";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011100011";
   IN2_i <= "00011011110100101";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000111110010";
   IN2_i <= "01010100101101000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110110001111";
   IN2_i <= "01110110100111000";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101000011010";
   IN2_i <= "01000100110001101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100010001";
   IN2_i <= "00000111011001011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010110101111";
   IN2_i <= "00100000101010011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010000";
   IN2_i <= "00101001001010011";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011000100";
   IN2_i <= "01010111001101111";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001000010";
   IN2_i <= "00011100110100111";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011011010";
   IN2_i <= "00111101011000011";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011011";
   IN2_i <= "01111100111100111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001001110000";
   IN2_i <= "00101101011101001";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110100000010";
   IN2_i <= "01000001010010100";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110111011111";
   IN2_i <= "01100010000100100";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010101000";
   IN2_i <= "00001110001000101";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111111101";
   IN2_i <= "00100011111100010";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011010111000";
   IN2_i <= "01111000000100101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100010111";
   IN2_i <= "01010111000011010";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010011001000";
   IN2_i <= "00011101010010001";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011000111010";
   IN2_i <= "01000010000100101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111111111";
   IN2_i <= "00011111111010010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011110100";
   IN2_i <= "01111101010110001";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110010010001";
   IN2_i <= "01010100111101011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001111100";
   IN2_i <= "01010110010111010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001010101101";
   IN2_i <= "01001011010010011";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100110111111";
   IN2_i <= "01000100110110100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100110100111";
   IN2_i <= "01100111000011000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011101101";
   IN2_i <= "01000101111010110";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100011011000";
   IN2_i <= "01100010100001100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001001100100";
   IN2_i <= "01110101100001011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001010010";
   IN2_i <= "00001110100000101";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000111000001";
   IN2_i <= "01100000011100101";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100111110111";
   IN2_i <= "00001100000011100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100100001";
   IN2_i <= "01010001111101100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100111111";
   IN2_i <= "00101100110001100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010001011110";
   IN2_i <= "00000110100001010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110111111";
   IN2_i <= "00010101101000111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101001101100";
   IN2_i <= "00001111000011101";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100100001110";
   IN2_i <= "00011111011000110";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001100010100";
   IN2_i <= "00000000011100010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000110000";
   IN2_i <= "00010110111010100";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110011010010";
   IN2_i <= "00001101111000101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010110001101";
   IN2_i <= "00101001001011101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100010100111";
   IN2_i <= "01111101001110011";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001001011";
   IN2_i <= "00100011001001000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000100000";
   IN2_i <= "01100110100010011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111000101";
   IN2_i <= "00000001011110100";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000101001110";
   IN2_i <= "00101110000100000";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011010110";
   IN2_i <= "00001101011111111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101001101100";
   IN2_i <= "00001111000001111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110000000100";
   IN2_i <= "00100110111001111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001010110110";
   IN2_i <= "00101000101101000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010100101100";
   IN2_i <= "01010101101111101";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011101011";
   IN2_i <= "00000101001101010";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000110011";
   IN2_i <= "01010110000111011";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011011100110";
   IN2_i <= "01101010000000000";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001001110";
   IN2_i <= "01100101110001101";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010110110100";
   IN2_i <= "00011000111010010";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100000110100";
   IN2_i <= "01100110100111001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011010010";
   IN2_i <= "01011110101111100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001111010000";
   IN2_i <= "01100001100010010";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000100110";
   IN2_i <= "01001000100100100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011001000000";
   IN2_i <= "00100100100100110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110111101100";
   IN2_i <= "00011100011101000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010101001000";
   IN2_i <= "01011010100111101";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000100011";
   IN2_i <= "00010100100111100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110010000";
   IN2_i <= "01111111111001010";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100001010001";
   IN2_i <= "01000011000000111";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011000111";
   IN2_i <= "01001100110000001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100000010";
   IN2_i <= "01011111100111110";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111010110101";
   IN2_i <= "01111000110100011";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001001011";
   IN2_i <= "01100101100110110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111011010";
   IN2_i <= "00011100010111100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110011010101";
   IN2_i <= "00000110000110101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111111010";
   IN2_i <= "00000111000100010";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101001000";
   IN2_i <= "00100100101111110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101011000110";
   IN2_i <= "01110000000110011";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011100010111";
   IN2_i <= "01010110001011010";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010100011100";
   IN2_i <= "01010001000111011";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110010110";
   IN2_i <= "01001101001000000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011011111010";
   IN2_i <= "01001010101010110";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111110010101";
   IN2_i <= "00010110000000010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100111111";
   IN2_i <= "01011000000011100";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001101000001";
   IN2_i <= "00010110100111001";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010001110000";
   IN2_i <= "00101111101111111";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000100101111";
   IN2_i <= "00011011000111010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111100010";
   IN2_i <= "01110010100111010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010101101";
   IN2_i <= "01111011110011000";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110100000101";
   IN2_i <= "00011111011000010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101010100";
   IN2_i <= "01110000000111101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101100111101";
   IN2_i <= "01110111001001111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110100001111";
   IN2_i <= "01111001110100101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011011100";
   IN2_i <= "01011001001101110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110001011001";
   IN2_i <= "00000111111010111";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100110000111";
   IN2_i <= "01101010100001100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001000011101";
   IN2_i <= "01000110101011110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011100111010";
   IN2_i <= "01100110111001000";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100111000110";
   IN2_i <= "00001011100111111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111100000";
   IN2_i <= "01101101011011011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101001101";
   IN2_i <= "01111101011111111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100110111";
   IN2_i <= "01000001001101110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110110010000";
   IN2_i <= "01010001110000011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011011001011";
   IN2_i <= "00100111101000101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111000110";
   IN2_i <= "01010100110011001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010101011";
   IN2_i <= "01011101010111110";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011111100";
   IN2_i <= "01111001000101111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111100100001";
   IN2_i <= "01111101001011000";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110000000001";
   IN2_i <= "01101000010001111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001110101111";
   IN2_i <= "00011111001101101";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111001000";
   IN2_i <= "00000011011110100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000000100011";
   IN2_i <= "00110101011111000";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101101110010";
   IN2_i <= "01000111101010011";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001100010";
   IN2_i <= "00110011110101001";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010100010110";
   IN2_i <= "00010010110101000";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111101101100";
   IN2_i <= "01010111001100010";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000001000";
   IN2_i <= "00000110011110101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010011000";
   IN2_i <= "00110111011101110";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111010100101";
   IN2_i <= "00011100111011111";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111000010";
   IN2_i <= "00110101100010111";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001001101100";
   IN2_i <= "01101101010110101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100001111";
   IN2_i <= "00110111001111110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000101001001";
   IN2_i <= "01110111110011110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000110011";
   IN2_i <= "00010000001011110";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010100111";
   IN2_i <= "01101010001100110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101111001011";
   IN2_i <= "00111101111000010";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010111011";
   IN2_i <= "00110000111110100";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111101011";
   IN2_i <= "01010100101101111";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101100001";
   IN2_i <= "00000110101101010";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010010011000";
   IN2_i <= "00010010000000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110111011011";
   IN2_i <= "00100000100001100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011110000101";
   IN2_i <= "01111001011110101";
   IN3_i <= "0100001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111001000101";
   IN2_i <= "00010000001101101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011110010";
   IN2_i <= "00010011001110100";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101110111111";
   IN2_i <= "00011100100011010";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111001111010";
   IN2_i <= "00110010011010000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110111010100";
   IN2_i <= "00010100111000101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101000111";
   IN2_i <= "00000010111111001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011010000010";
   IN2_i <= "01000111110010000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110111011";
   IN2_i <= "00011010000010011";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001000011";
   IN2_i <= "00110011100100111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010001001";
   IN2_i <= "00001000011101001";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001000010100";
   IN2_i <= "00011111100011101";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011000001";
   IN2_i <= "00000000011000001";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000101011011";
   IN2_i <= "01100010100101000";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101010101000";
   IN2_i <= "01100100100110111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111110011000";
   IN2_i <= "01000101110100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101111";
   IN2_i <= "01000000100110111";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010010100";
   IN2_i <= "01000000000010111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011001111000";
   IN2_i <= "00111000101110000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001100101";
   IN2_i <= "00001101100110011";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010111111001011";
   IN2_i <= "00011001011110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101001100011";
   IN2_i <= "01100111101110010";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100101010110";
   IN2_i <= "00011110000110000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011110110001";
   IN2_i <= "00111100001000000";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100100011010";
   IN2_i <= "00000110001001010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010110010101";
   IN2_i <= "01101000011011100";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111101000010";
   IN2_i <= "01100100010111000";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101111100";
   IN2_i <= "00010000101100001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011011010";
   IN2_i <= "01001010000001101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001010010100010";
   IN2_i <= "00000011111110100";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011100011000";
   IN2_i <= "01100110000010010";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111011111110";
   IN2_i <= "00001000000001001";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000100111";
   IN2_i <= "01010000110111110";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000011010";
   IN2_i <= "00100111111010010";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110111010";
   IN2_i <= "00100100000010010";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010111111";
   IN2_i <= "01000010000100111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110101110000";
   IN2_i <= "01011111101001100";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110000011110";
   IN2_i <= "00010000110100010";
   IN3_i <= "0001110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010000010";
   IN2_i <= "01111000110110101";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100000010110";
   IN2_i <= "00101010010111011";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000010000101";
   IN2_i <= "01000111010101011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110000000111";
   IN2_i <= "01111100010111100";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101000101011";
   IN2_i <= "00000000101011100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001100100111";
   IN2_i <= "00100110010011101";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001111110";
   IN2_i <= "00111001111110000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101100010100";
   IN2_i <= "01001011011010101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110110110011";
   IN2_i <= "01101000010111101";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101000011000";
   IN2_i <= "00111001011000011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101000101101";
   IN2_i <= "00000101000100011";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011001000";
   IN2_i <= "00111101011001111";
   IN3_i <= "0010001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000110010001";
   IN2_i <= "01000100011000010";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110010010101";
   IN2_i <= "00100110011111110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011101010000";
   IN2_i <= "01111101000111001";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101110011111";
   IN2_i <= "01010111100110000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100111101001";
   IN2_i <= "01001100011011011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011111111000";
   IN2_i <= "01110100000001110";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101111110100";
   IN2_i <= "01010011010011011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011101001";
   IN2_i <= "00010000111111111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001011100001";
   IN2_i <= "01111110111100001";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011010111";
   IN2_i <= "01000101100110111";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000111111";
   IN2_i <= "01000011100100100";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111001000100";
   IN2_i <= "01000011011101100";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011001010";
   IN2_i <= "01011101011111000";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100101101001";
   IN2_i <= "00101100001111110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101000100";
   IN2_i <= "01110101111110110";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001111111";
   IN2_i <= "01011100110000101";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000111101111";
   IN2_i <= "00101110101100101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100001010010";
   IN2_i <= "00000101111000000";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100000110100";
   IN2_i <= "00101011000001000";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110001111";
   IN2_i <= "00010101100101111";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000001000";
   IN2_i <= "00000111101100101";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101000100101";
   IN2_i <= "01100011110010011";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000000000";
   IN2_i <= "01011010110010000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011010010101";
   IN2_i <= "01110100001001111";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111101110010";
   IN2_i <= "00011101101101111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111001000000";
   IN2_i <= "01011001111101001";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110001011001";
   IN2_i <= "00100001001100110";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011001010111000";
   IN2_i <= "01000000100011011";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001100011010";
   IN2_i <= "00001000101100100";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101010001111";
   IN2_i <= "00110101001101100";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110010111111";
   IN2_i <= "01000010000110011";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010011100";
   IN2_i <= "01001000100111000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111000000000";
   IN2_i <= "01100001001111010";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000010001110";
   IN2_i <= "01101010101110011";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001001100111";
   IN2_i <= "00100111001101000";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101010101001";
   IN2_i <= "01101011011110000";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110001001";
   IN2_i <= "00010001001010100";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110101111111";
   IN2_i <= "00001100110011011";
   IN3_i <= "0011111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011100111100";
   IN2_i <= "01101101101110000";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100101110011";
   IN2_i <= "01110100001100110";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101000001110";
   IN2_i <= "01111000100001111";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110100110110";
   IN2_i <= "00100111100101111";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000001001010";
   IN2_i <= "01101100101111110";
   IN3_i <= "0110000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000001001011";
   IN2_i <= "01110100000100001";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000000000011";
   IN2_i <= "01100110010001110";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000110010111001";
   IN2_i <= "01100000010011000";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110100011001";
   IN2_i <= "01111001111011100";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000110001110";
   IN2_i <= "00100111100111100";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011011100100";
   IN2_i <= "01100101100010010";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100110101011";
   IN2_i <= "00001100011001111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001011110101";
   IN2_i <= "00110111000110001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001010111";
   IN2_i <= "01101011011010001";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001001000";
   IN2_i <= "01001001110100110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001110110001";
   IN2_i <= "00011110011001101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000010010000";
   IN2_i <= "01010000001011110";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011000110001";
   IN2_i <= "01101100111000110";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000000011100";
   IN2_i <= "01110100001011010";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011010101101";
   IN2_i <= "01100110110000101";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010101100111";
   IN2_i <= "00110000100110010";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000011001111";
   IN2_i <= "01111100101011011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001111100011";
   IN2_i <= "00001001110101110";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101000100";
   IN2_i <= "01101101001000111";
   IN3_i <= "0110111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110010110";
   IN2_i <= "01111100101110011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111111110";
   IN2_i <= "01110000010000010";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111111011110";
   IN2_i <= "01000111101011000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111010011101";
   IN2_i <= "01100010111010100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110111011";
   IN2_i <= "00111000000010011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000010001";
   IN2_i <= "01000011100011011";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110010011";
   IN2_i <= "01011000010101110";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011011111011";
   IN2_i <= "01001110101100110";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011110111010";
   IN2_i <= "00001101100000001";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001101100101";
   IN2_i <= "01101110100100101";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000011001";
   IN2_i <= "01001110001011111";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100001010";
   IN2_i <= "01000111010000101";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110110001100";
   IN2_i <= "00010000000010001";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010001110";
   IN2_i <= "01000111001101011";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101101010000";
   IN2_i <= "01001110111010001";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101001110110";
   IN2_i <= "01101111101000111";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011101010000";
   IN2_i <= "01101100111111001";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001011100110";
   IN2_i <= "00010101100101010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100100010100";
   IN2_i <= "01101111100001101";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001011000010";
   IN2_i <= "01001101101111001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101110011100010";
   IN2_i <= "01101110000010011";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010011000001001";
   IN2_i <= "01101010101111001";
   IN3_i <= "0011011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111110101110";
   IN2_i <= "01001001110001010";
   IN3_i <= "0010010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111111011000";
   IN2_i <= "01011111110110101";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100110101000";
   IN2_i <= "00010000101010101";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011001000";
   IN2_i <= "01110111001001101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101101000001";
   IN2_i <= "00111111011010011";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011010011";
   IN2_i <= "01101100100010101";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111110101011000";
   IN2_i <= "00110101101111110";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010110001";
   IN2_i <= "01111001111001000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000111000011";
   IN2_i <= "01000101010100101";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000000001";
   IN2_i <= "01111000111011000";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001111111011";
   IN2_i <= "00111110110100101";
   IN3_i <= "0111101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100011111";
   IN2_i <= "01010011111000111";
   IN3_i <= "0100010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001100110101";
   IN2_i <= "01001110001001100";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001101100";
   IN2_i <= "01001000011010000";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101101110";
   IN2_i <= "00101010111010110";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100010111";
   IN2_i <= "00000110010010110";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000110100011";
   IN2_i <= "00110110010010101";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100011011000";
   IN2_i <= "00110101001011011";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100011000111100";
   IN2_i <= "01001011000101000";
   IN3_i <= "0101000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101011110";
   IN2_i <= "00010010101011001";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111100001";
   IN2_i <= "01010000110010001";
   IN3_i <= "0000110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001010000111";
   IN2_i <= "00010101000010101";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111110111100";
   IN2_i <= "01101010010000111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000001111011";
   IN2_i <= "00110011110000101";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101100100011";
   IN2_i <= "01000101101000011";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000001010";
   IN2_i <= "00001011001001101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000011111";
   IN2_i <= "00010100000110010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110001001101";
   IN2_i <= "00101111010000100";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011110010010";
   IN2_i <= "00100101011011010";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001011001000";
   IN2_i <= "00000001100111010";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101011001011000";
   IN2_i <= "00000101111111001";
   IN3_i <= "0001000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000101110001";
   IN2_i <= "01100110111100110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000110010";
   IN2_i <= "01011010010111010";
   IN3_i <= "0110010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000000111111";
   IN2_i <= "01010110111001011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111100010101";
   IN2_i <= "01000111011111101";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111110101";
   IN2_i <= "01010101010011010";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110101101010";
   IN2_i <= "00111000100110010";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110101010010110";
   IN2_i <= "01000010011100000";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001110011100";
   IN2_i <= "01001010111011111";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001010101101";
   IN2_i <= "01010110101010111";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000001100011";
   IN2_i <= "01110010101011000";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100010000010";
   IN2_i <= "00010001010101001";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010101100";
   IN2_i <= "01001101001110101";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010111000011";
   IN2_i <= "01101100110100001";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000011011";
   IN2_i <= "01011110010111101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001110010110011";
   IN2_i <= "00110101010011111";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010010100010";
   IN2_i <= "00000011011000111";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000111111010";
   IN2_i <= "00010100111110011";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000111001111";
   IN2_i <= "00100101001110100";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000011101110";
   IN2_i <= "00011011000000000";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010110111010111";
   IN2_i <= "01001110001111001";
   IN3_i <= "0011101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010000111000011";
   IN2_i <= "01111011111011110";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000100110";
   IN2_i <= "00000011101001101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101000011110";
   IN2_i <= "00100101000001110";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101101100011101";
   IN2_i <= "01110011111100110";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100001100111";
   IN2_i <= "00110110101011101";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110110010001";
   IN2_i <= "01010101001110100";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010011111110";
   IN2_i <= "01000001011011100";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110100011011000";
   IN2_i <= "00110000111101111";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111010111011101";
   IN2_i <= "01101100110010000";
   IN3_i <= "0010011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001011100110000";
   IN2_i <= "01110011101011001";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011010011001";
   IN2_i <= "00110111011111101";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010001111100";
   IN2_i <= "01101010000101000";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011000111";
   IN2_i <= "01010011111111001";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011111111101111";
   IN2_i <= "01110100001100100";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101111101011";
   IN2_i <= "01011011011101001";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010100011001";
   IN2_i <= "01100001110100100";
   IN3_i <= "0111001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001011001110";
   IN2_i <= "00110011110101001";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000100100001";
   IN2_i <= "01010011100001101";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100010000100";
   IN2_i <= "01100001000001001";
   IN3_i <= "0011010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000100011010010";
   IN2_i <= "01000000110110101";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110111100111010";
   IN2_i <= "01100011011000101";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001001011010100";
   IN2_i <= "00100101011101000";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000010010001";
   IN2_i <= "00110101111111000";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010101100101011";
   IN2_i <= "01011101011001011";
   IN3_i <= "0000011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011011000011";
   IN2_i <= "00000011100011100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101010100100001";
   IN2_i <= "00100111101110101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010010000001001";
   IN2_i <= "01100011000100001";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010011100110";
   IN2_i <= "00000111001011100";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010001110010";
   IN2_i <= "00000100011001000";
   IN3_i <= "0001011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100011100";
   IN2_i <= "01001001011001100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110000100101111";
   IN2_i <= "01111100001010011";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001010100110";
   IN2_i <= "00011010111000101";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100111100110";
   IN2_i <= "01100100111100111";
   IN3_i <= "0010000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100111110101";
   IN2_i <= "01001000000100011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110011111";
   IN2_i <= "00010100101010100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111000011111";
   IN2_i <= "00100111001111000";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100000100011100";
   IN2_i <= "01011000110110111";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000010000110011";
   IN2_i <= "00101001110110110";
   IN3_i <= "0010101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011011000010";
   IN2_i <= "01101100001110101";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001100101011";
   IN2_i <= "01111100111011111";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111000101111111";
   IN2_i <= "00001101010110010";
   IN3_i <= "0000111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100100010000111";
   IN2_i <= "00001001100001101";
   IN3_i <= "0110011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101001000111001";
   IN2_i <= "01111000111101100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000100111000";
   IN2_i <= "01011001010001000";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000000000010101";
   IN2_i <= "00100101101010110";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110011000100001";
   IN2_i <= "00000111111001011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010110101101";
   IN2_i <= "00111100100111000";
   IN3_i <= "0101001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010011101111";
   IN2_i <= "01101111100110011";
   IN3_i <= "0000001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000111111111001";
   IN2_i <= "01101011110001111";
   IN3_i <= "0001001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011011110011000";
   IN2_i <= "00010001011110011";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000001011011";
   IN2_i <= "01001000000100111";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010001000000001";
   IN2_i <= "00101011101010011";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110110101011111";
   IN2_i <= "00000001010111100";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001100100100";
   IN2_i <= "01010111111001011";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010111011000";
   IN2_i <= "00001010001110101";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010000001101";
   IN2_i <= "01110000010011101";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000000100100";
   IN2_i <= "01111100101110111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011000010000000";
   IN2_i <= "01001011011010001";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110001111110110";
   IN2_i <= "00000111110101100";
   IN3_i <= "0101110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001010101";
   IN2_i <= "01111111000000010";
   IN3_i <= "0000100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011100111111010";
   IN2_i <= "00101000110011111";
   IN3_i <= "0111111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111000100101";
   IN2_i <= "00110101000101011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100010100110";
   IN2_i <= "01000101011001101";
   IN3_i <= "0011001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100111011110100";
   IN2_i <= "01100110100101110";
   IN3_i <= "0011100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0110010010010000";
   IN2_i <= "01011110011010100";
   IN3_i <= "0001010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111101011110010";
   IN2_i <= "01000101110011001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011110010010100";
   IN2_i <= "01000000110101101";
   IN3_i <= "0011000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011010010011";
   IN2_i <= "01010110111100101";
   IN3_i <= "0001111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110001001000";
   IN2_i <= "00100110000110001";
   IN3_i <= "0101010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100101011010";
   IN2_i <= "00110000110100000";
   IN3_i <= "0010110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101010111010";
   IN2_i <= "00000010001001100";
   IN3_i <= "0101101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000001010011010";
   IN2_i <= "00000100000100100";
   IN3_i <= "0000010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111111101001111";
   IN2_i <= "00110011010110110";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010111011011";
   IN2_i <= "00101011011111010";
   IN3_i <= "0100110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000101110101110";
   IN2_i <= "01101001111111001";
   IN3_i <= "0111100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010100010100";
   IN2_i <= "01110010100100010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100100101111";
   IN2_i <= "00001001111110010";
   IN3_i <= "0010100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101011001100";
   IN2_i <= "01101111000101011";
   IN3_i <= "0111000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0000011101010100";
   IN2_i <= "01111111001011110";
   IN3_i <= "0110001";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001100110100000";
   IN2_i <= "00110101101000101";
   IN3_i <= "0110100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111101111001";
   IN2_i <= "01111100110111000";
   IN3_i <= "0101100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100010011110100";
   IN2_i <= "01110011110001110";
   IN3_i <= "0110110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001110011";
   IN2_i <= "01001011011110111";
   IN3_i <= "0100000";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001111010100110";
   IN2_i <= "01010111011000110";
   IN3_i <= "0100100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011010101100001";
   IN2_i <= "00000010111101010";
   IN3_i <= "0111010";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001101101001110";
   IN2_i <= "00111100110110111";
   IN3_i <= "0111011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100110011011111";
   IN2_i <= "01010000000111000";
   IN3_i <= "0001101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101000011001110";
   IN2_i <= "01011111010111100";
   IN3_i <= "0100101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0010100001000010";
   IN2_i <= "00100100111000111";
   IN3_i <= "0010111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100001110100110";
   IN2_i <= "00111000011000100";
   IN3_i <= "0111110";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101111011011101";
   IN2_i <= "01101100101000100";
   IN3_i <= "0001100";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111011111111010";
   IN2_i <= "00110001100001011";
   IN3_i <= "0000101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0101100001010101";
   IN2_i <= "00111100101001010";
   IN3_i <= "0101111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111100011001101";
   IN2_i <= "01011010011100011";
   IN3_i <= "0110101";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0001000101011010";
   IN2_i <= "01100111000111010";
   IN3_i <= "0100011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0111001101010000";
   IN2_i <= "01001100011001111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0100101001000100";
   IN2_i <= "00110101110111111";
   IN3_i <= "0101011";
   SEL1_i <= '1';
   wait for 1 ns;

   IN1_i <= "0011101000100010";
   IN2_i <= "01111111101110111";
   IN3_i <= "0100111";
   SEL1_i <= '1';
   wait for 1 ns;

wait; 

end process; 

end test;